`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PPW701Ppq73bxe3/y7KZEx571fPBQyMSRVmxs8QhJrJEMPP+NW7otihnCjq6cBv
jYYgILPc4xG/VekWh6oezU7rE60yTqlUHz+zHTgMHHygwXsl3kfrSliuxBW07Jpt
g/vWLDuw/Je3bs5ln8v4oTPnKvyk6MD/4PK7SoZJ/Ckrrpv+ZwswEdx/A4zrwmT0
03puu4jiR9mLZ0nTvhdfmJwM+oH0GfzW2h5BPQwEfjhS5CCMl75S0z5uxOvYYotL
xaN6kToxvHjEdB+hjF4jYk/c3ruvNuA2qUGiuIaftU0FJkb74K18D/CHIkCHTHD0
IGDPZenx3AVvA1CcCLHyQ8+AkGaBginBpucKadmXi9YFJLPGKoujHY0VlNRnod/n
1eCCUo3/V+3EUFsRDl/W+eoml4nKnLr7LFYma8XH48geoxcYxhngS7U4COZN9cL0
drTsz4jriwV3KrkQfyLckyIRaolNAJl2S8CSXYzjEGpWJTZpX1zu2TWA2IeUBuiF
2gnW4S07dxDHOx0ra33s9Xv4LFH7tAk4i/JzLll7t6bK7OkM38YsDW9x3UCmtzWG
XHUew4YeLbC7uGNCc1g2zjSTkTqSlTEThZgA9CScomBXVqCArw0yyDaYITanLxmr
7fIW2dnnNEOoszTeFehOXnNZZsv4S34THfWpKEvP5thBSLYJIc7cY4UpssxKisJg
c6YRJWlpk0HcrpJmDvfZbdCaDpospKtdNQv2l+7jeND4AzmRfXBEvXmhVkm2iVxJ
LV9lsInownsP922UPYi1AgVktqfCM9lih425QiFiHtpTSgHVNMvsilOOe3AQWcQC
i/dZr9FsLkI7gc7ezcy7MBr/pOD+r8GnRWMocFO9abXKbAQ/MZJ7uGq4mq1NqFMl
nsfRSWZzA+SsMiiq9bzHQZwM8ZRd5jfhvxg7Upqa7Bl/ytyudiE4OqzON0xwfjjx
/fxMweXjJVd/qygqc99dCZvRAouCGb7kVPYMJuoxcfjiTbElY+l4hgroRXC6+VLG
Tltcv0+BZZ7K4pgKeBTQia3BUr1dTC3RwnTPPjfELri0zOvCUudvk31gvhqlfsz7
RM+wVHNIb5Q+fCeKbkk+9RTQ4XXVwFP75Pqr78XN0F93qEGB15/nd3lqJim1sLuy
zr52O6nOfVHcHxPZIaUs7vhhVAmjqpYEqjxhMQRiudy5l2xRMRaONg8+CsS1snua
VTGbWAMUykJuyHpywSVmu/pOGQIiKj1gNYtjgWPyiJMbTyON8EcFsvp2Mv5FPk5z
/QKUgmSxgct0vm3nHu+Z6tf6i5ObmXDgR7GxCySIXMPTBQzI2h3hPbQREF8uDgjn
fCyM3Ia4SEs+QAdoi0s+F+Q0hYeJETu1U5nH62K8F/QX2lTmJ4DgPKlvZZWHd/iP
+oreFLniIC30+qdIYGKSQVWAl6xZqsEQylcZ0eLaABNvNLXKHqWubCZhhL0XRkZg
Ec9I0CxyMHeqYTF0fOF/awCJNToijFtCs78U9z0G8EtSW8HkU935SfVHzPDrW63O
tckEH7RQc3h2hEPxX5E3FVeKwfAjBQEfY5my2mL28G3pbII44VaAsAW28fDVleha
l4FAWuid9atSwuCqMiZWv3bHaZ51nIGgmwqDFPkagjRfRj9Hab0nQqcUwyg7Wqde
aR3kjT7dwRDprzk2c7g5arn7/kID5F3XuD6C6M/zUqOA38VoFWY9Afy3AJq1uZI3
69ChUWDiP6cum8XNXVmD94g5peNozlAUdjnq6f3GRK0XUsgyjV5fCviOJI6CCTDW
MO7COyrnRs0imvSZLoDH7hvwa4/crY7qjI/W7iXVISjU+84jh/dwu8YpvfaKSPnd
iTcFGJNdjaynOIcT4h4hsg==
`protect END_PROTECTED
