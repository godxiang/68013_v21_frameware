`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEAfETp0m/nO4QiagPnCHnfrziuWFxuSYvHoooSwE4d30uZO2rMfIc58jCCBdIqd
/XIF0g46tIqMa+heItU/+7RftUr0ENguvFtR6B6WgcgeA4u+ZUCqdEb2g5ERuBQe
93m0EY4j8D8DAKj/SEDxxhxITCXYSGlMldjbQusgdOPc6Mx3mxx2SDkDz1DwJOa9
5iuzXDhXjbu0LtrfracPB/m9qhQ9u8tBTeMcrz6RYEH8sB2bTSuEoKgBD4fL4Rdh
GWFPxl6RqwrjQ0ZvPn7VORtptCYgF5ngFVga5ZVTQHGCuS5oDFWEAu8QxeVp9MoW
9qRqL5GW8YwSUhRrzDUAI8tRCpxZVCSEjpNFHcJJP8HU5szGWDaC4PomJ5GgkAAT
C5S1bxkud+EC1dEGcjwVyhc5KavZ5SNzb0cnnhMT+2utIlU6oZxkM8FoIPwAiFWR
peTDS1QEw8WvoVg+jMNPor8azi+qYXkuaPGykl4L1CkgxB5+novwM1tZnP8bi+sC
xNM5Ff9ZBTkmlf3znGafFI0BRCUEx81VPboNvWI4OLc1kOC/wPCEssRJgOPztrGx
pnL6blE3N+5oaiky/mhPDPond5jaLBjw4o5QoX/w7NABivFVBrJOMebTM5ldZue1
xDGoMumE2ngL9b1Qv/vLoo19zzly6MvqRH5GBi+S+ZdCHOQcz1ca+wuBliCxiXRw
m6fz4RWc4Q4R1idIc/j7ifiNqQ/bUPDNZHWcRtxdK0sIjsxSwZ9prI5w0/68v31L
J7PgSTcnAsGFSNnb9J2logR96MNc/35MSQCcSPe0u92IAbf1cOn0bzLreN/3Kx9A
4SaYKqJLj/CVFWySbvGp9KikMGQJbDLacR7eQoyndS4m/8iyBdaJPoRasWRTwyrk
n7vu11K7oITFPje3sSUoW7h94O32ax7FMzi6bh40f2yJL9WnprJ/dPfc89KHWLSg
Zo+6CvSkEr0vqSQdykHs4PL7UGWSDkWduCrm1r2wZpFCwEx13XtpX4ZvrM+aZpvQ
GvQxJ5FUhTC9edutWxWMaInaKZS3oX82aDhYk4xl0kRY/2oCA+mQK4Xt1Y/KqxAT
vWCv5M2/J+3pImDmbTzytwDY1N3QCt/p2DDjvf8wLryncdSIibSeXZc0w6p5YIVs
p+nOW1dkMVAjmqe3S9QXULVt1Mt4N8uHYrE4isWp7Q/3T2KzqNbeJynZtNyQpuTN
yIriqdaPxJNbP6FOYsEskEPOunpi/HJVxgWpRF75rJhzSIc6CLFdwmoC7YElR3V5
Zo+tI4GTZeqmGi80IiGGJ1VOw16yWWE15Iif9zki+YnzctQSGXZWbGRaRdQobf9s
RB+VCKuL9JF3R+G4Ypq9KhS0A6yJgmUhgKrJUq/TUtzBr1SvzgeGeHd44IpA+lDL
WeOX02iGlGF7uRS9lN5vxWmX+QMgzkqm5d0AR5DUX/jIR2tV0mF99WzSoKQFPv3n
59zC59DiI/ZU48KU1a65YahldNI+RrIdVAp8CAM05c34cZVD4S5cVLjVlOQ/iUEA
k26qB8/Kkrg/GJQXBgRFZdm60jS3//RZa3qAQkVFvJBzjfNPct2lwZdKioygjxmY
s6CsZeDLe1llAhdlsmDNmTWK5h6cgXeeQFEeAK5WzQ0dIrWPGRx5GzJepRY3mpbK
qyc48QhhAoHpGSA+9s+x0TmX26iMpGxU2zn0hh+jB1znf5Auej38PiC1sl3O3sOZ
5iUz5Tg9ynURrwOCCFtm4spCIaP18TGqh6voVPtHmNT/ranAMGfn9/ERPyJnano0
e1JHFdE7RJlvc2pyO+D2hmknEdSUwN757LEVJwQ61jO03inEfoFKtu3IYeOQfsgb
0qcj62XWSPnXX7KN1vt9JIFH5yG6qi5mAgw81tFDg9IaOuoXPNWpQbp6qds5EbFN
PTZrjHrbe5zZBYyXThoneIBNwCtSb68tiu6GRBi4In46QRjLMRvz+0Sa/AsKHTfn
0Db6YO/bkgKhtJtrABH438aJdy21f0zJB5iFhJXzc1spy0wdxX7Z43+KjZlCXVo7
1wQaQcYYbVWjyNrZ9dCLEP+pUFt1gN6vVEaHauxq8daJLVSrRSCWF7SnBDLlOz10
4lT+Yaal1YR0hEtCJG4DFzV6TJwvQNodUIwdLX09y0H9+IZcHgnocy7K5KWEVh2b
Fi+tBu4HYiKzOgjyKos5tuSh1bii13gIUFE/0kBexbrmtV45acPkvdloipMLMdzh
MjzjGLkrh17KQVPjmDHUF7wH6BivHs9d0pKRYoOVZ9MdFNMsyQaboTB607+9h/1d
vBFu5SQ2KyUJ4Zawv+ryQ5DPHSi70kCxUpvL8OGgNREM43dRRHT20yXrJxCsjunH
zas6HNCs2LFIIUVpOawytEyJxrDffcHFtYWfU1LVt63ApBXKcsgYBFiLxSQuDRjR
EpGjgn/9mZKVVFAlHBUoW8a42dY+3s/e2ug6zfKqJEiCYbIqEN35JY8CoGem0+jD
66BO4M0BZ70sXvQVWSNburpJ+SSmHghCew8qAQHQrtrCZbq24QCWutbETmrC7as4
tyaZ6kpnfRAR2O0rvffGL+/MiFjr3ciUhfKnTyqYLuUnYPowKjiV3DFcqgqwPSR3
J9pOA+J2TPpyyBdbmMOii4HUXT8cGxWToFWA4DsM1OZ4JpasaMAiRPKnnfcpKkWx
5g6r50taFokPR7zuDj/qaO5omSVcTob0jwMbgzJOpD3PboRLn0O+vhuUcmGNAhK0
7FJVV8mGAJJMfjEWtW7bOvU7RY+rVoZTZpMQjV4Wesg/HhOYLL6QbjWko4XABSym
2d3FKuwX70FL+uLFyEBZtZtyHtEgak9b+fmYZGOfXsDu0ayDMP3yCJUo5QExiCqZ
2tebhS01oVhCNhS5MKiizGZ5L6VY1RIu+QXTIpRe0xCsPpaKsCo6gO6JQKrQyLDk
egB+POIOyE+kKovMru7vE6y1fsvFGgPZ/qDIa5V0nbF+lb/GRpajQ9G0iK7RwuLb
QE8uQt4JvssyQbLkf90uiBPqEUtsqDLI7Wj117W1bvlDoe4uXXsNYtdyC6h9SjTh
6d5QPpXJUOhn6dzKVgpYc4KNyMO5py3IIKhgFCQr/RrM3yuMoO4MDS2f8vAj8NbR
VM+HGlS2oDTmPDQOhMPoTEOyth/+SlDUxxcveJU7svFoDVjf9U2k6MvoMX2qfjKn
bFZDf9kNQSRTfGse8ZKWMCYLj6QHi9dlj4NtK46BAgsYCMAFeOV1viNk4tzokcaE
Kn2V1WXVD5A7q/NkFdp1AeYRCdI1h7KkjJAOxUThxnAoyybYSQWoCa7i0R13k6Al
SReOwalVTUxvouiXX+pXkB+h1F30b9f3xHIjRuUnJdqHizfFARlpBu17O/LOvYeg
33Sy+zv0U0MkrWW06ZHXkOrELaPDBzQp+zsA0S7KFB5O7abUtJo4ZncQXCT93zG3
PfQB7198aRtcfI4PGabeOwwEjkZS3Pjmp1d9WBcH0JKEINRYxhFXRiIMitDSv/Gt
72Vn6EeKuANbqNOM1DeS+JnP2ZAgRNqT1oC0Ce4dahyrO0xS5WXGguP+IHeFeSh6
eOG51z62jmFtfpyLfdeBcZ345T4UBjgbobI2WtEu4ehQtj4FT+hLUjO3kvffqD2p
/ILfHVdErl6kyNr+t8q62v8kZGhN35hoFmvpHmZuVyZzAIk1PJ8iePWIib+uR7b5
172hqQDSDdAT+0/ghPIlwnkqsLplHkFhzDwF++1RQj+/6ff7+/4/qZBLTEgR1XIW
n8tKBpGo6UAJmXHcNJF+4Znh5bE0mMbyQFLjYLXUtTdTwo/CcrkPuiSqKWLupZay
FJif2JforaQA0/ETMpUQP0MKKuOVw+DLwRlXfYahMlNxs8Cg6ZzYiqVpB+BN+WF7
mT+i4wI/Iu1iM3y08+fBHlRo7swxK7cOlUUdrlQDE17eiie1OX3wEejJYhnc5MAR
BvDCz33CoPhnVea5q6AtINYrdjMiNpuX69hKpPf6WpehQPIDnbQrXZ0gW+NU2Naj
76l4pCyMzZeUqSoZH4S1Dyl+MAnnwYdamehHBvgVKzOe+ZMl+V4pM2RHrGxoO/NL
PpOHUYTmHwSz/fqMhfYCpKbEOrZIz3bLbf1AoaX7F6edq5mVU8qLmljo4Eb/Achj
akl+D/847ZX6izdcqrg7aRvdX5jAQOrLm8Fc8emq07tBUtEJw83GJMiyqB6abqDS
ZYQlmVt+YbPtWcJgvRDg7uuMrojSseLombPIJEwrTOirr0qhmc/gKwkd86oZDuZw
IRdT6EiHOvW21OAryYMRJIGeYCPUpCP5fjLMHV9orm6M+SbKfc/C6IUmjgqNtSON
ia7EiNVfrOt2jp2+FJwzHyJccFMnPW6h260SOhFDOQY=
`protect END_PROTECTED
