`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3u6oWYZpiMxS45J5bIi0wyv2jx5odPyXJ12CCIvsEQ6kWISc+pBE80oZKcJwEwK
ZEYUZ7OywsyeMUiMbbbEM2GQ9PVVzXh07hrw6rLVfaxu0gse6/U4yWaOX7wNTcjC
w34+lyQ7QuVOiLH0Ui51T7gK+9sLsJzsnGqej+Xq1gtxwNnDtBVnNqI8wkqVx9Gf
p47mTka8dMRaD6xyoZDWMIls4xFKob/mPzzP1mEkwwVRH5ZsQxrCm33aqqSrG5F8
sgmB1vLdlYp499cpjhKm3rgDrgzC149FPU8TZG4fmlSF3Wm9JpFlrPTbkKseaVXJ
1ssppNgDGzvyAD8fKorEHMD6oYTQetyzR6jdztvlRVvAjlC2CqxLmVH7cgrIcrfq
`protect END_PROTECTED
