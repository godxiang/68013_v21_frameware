`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXwW0A3wzBcbpoaaHsdY8wSlv0bHw1QSvXYE0xn0wbXehG4a3V6DzZdXEWH1Xp/o
upThFImzruyNUZi/Y6zralRMUK54F8quCFy/dtdHNIm++mHobVjJNsfkDHEZqukc
u6S7invof4xZHk/kamAaFwwHkSEQ+vVcA1Tt4Yj8U0zDsB6SXt2YWpNHzuw5hG1a
Ww3tkq96AfRllxg/wDK73ngrEKo4FmZ1KC/aoZh2HVfri4N2tImlhJPnzKrKbH0o
OwVI09ZZ4Bv6w06FN4vqQfCN3L9fPEYpfLLgzCytyn1rDVSiOp7rA9Bc+5BZkjsu
4/0VcNhnyOyds632w77k2KIfCPwxbzHo0VpUYaj5B/6Ur5GimU75R2yg8N+yi3dL
uJ/+K+u+I43guaJwTDibrtwDA557IgIoBHeFdroRzdchvc200I/4sBgGoxnLfWrs
QV8QbqHatnxyhl8ADO03KtyX76LbrC4wlA3DLs9OT1burjnnbf/W+tQQIIhE2h/Z
mbZ6ZFB797qi0xU7RjY/LYTJa4ro+NcvGjLIrJ14aUMBS34kQtLHEQIfvKsGsyhi
lxnw1nAxcmntCxW6vNqo4HZHd3Uq89qmYb8sHjvn2TMg6mZHr/mNQ21505GT34hY
/ir33cXkN/mVRDNVCw2iZC3y2nnZcX1k3pnl5Qw7Q15ote3FFt8n4skEk//kdXXl
lhdhG/DWbWw8JBOJDjiOiM5oF6yZfL2reOiyON+h+cgJx1RBxfqVRfgX4DBoZ+LR
Rx4XhI7MKVodDK70EZFwFVuFGkuY/eRruJNKJZ1SVWdL1c3K+FrCkNwPtlMrWIwG
8zrODBScuGKu70YsXc0aJFQ51oKoIuQ73NYN+TRpXCPN8KoyxdVoS+IAkoh+J9Tv
fROXbbwxT46rkHBkEq4aXZzqcRxx08uu54Fm+4Nw6vKlX8gMf7ophYFkrsEitToH
HeU/FlYGyi+qLFYFLzlj6QEVscf5FRlsYeom3gRb5lVnSpFPNK66kUjvwLNpuyqT
jQxooQDcg9BcRVjKOr9Vhf95ZRI6DVauKVf0OhEIMK+20wVF60Asc7KPiBNNQmPr
`protect END_PROTECTED
