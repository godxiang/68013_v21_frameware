`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EcQdUbVlzpJJe851bzn+2ovKGV3i/T820hjTSbvzfriL/UKcVKypIKiVLadDSdxa
CTHUlRm8kDDA1FU84P7hM/zHRXaGtOQppZIk7ER5PW2GKhD91FO8zlhjnF0BiV4f
HjhjpNRnX8Ug2ETD7uUAwsuWs61Idj3jY8ipIVul3nrAEnjc9OcBQQ2bJlxgJGPD
`protect END_PROTECTED
