`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oj8SEFQsfb8+YAtqaSGv4LKQBxGjlQ92oaOYgdAKFOz9wYUjJAd89gkDXT4gB4qc
UTlHP7s5FG/5gT4tDgYg2X2hta0UUpXh73AJreLP2K1Ng39wYvHn8PwXnyQDVOR6
IdiAPZaRTZ1JprKeMQySL6BV64zhvb2EP9jzyqOMi1nMFwaR+I/FLqPTInjJeDWU
lbYjYpZYQi2I5h2VTBRsPMePacQaAqJjPM4Up8hZS2zbiftTfaOUY6TOdFXavZxJ
jxr/ewVLqMFQkxQSLXsZYZofk2ZUeq0me32Ce7AjVL0ZZuYFUSOTu5t0gT5OcFY9
DYCS621e6KXFw9FAITo4+1uhrtTAKPIA2pkiwUwD0KSqnuTv0JTQC2t5+fD+sBaE
eYz2zXvi/8tfrwYc6XYfqtksR5EIgQl0nQEAQ7OVkGbRMPgesJ4I1XYx7w54K/ao
9h/giPaeDj+fjR+Eq960//TtLt1ey+B/FlXm3KxL46WCZWdXc0BSSiabynbhPT6C
FOlfbyQqaVkAHuSeCWAIpE9YmoS2sj57hL4VxFDMOS2y0bC7cHpSv52utkjnYab9
1vK1R2n67YCOekMbIiOKAHUeY8oCTZjOteARBRagNFqFHu4XhgZG3YeiuOnh988W
v+R5rfWyrNP3oDmfC0x5mQYTkaigAJu+ZJa8HJVkqUq3LKGUclbK9xATChDDEwhV
g0RaoRzs6dSr6+YlIkDdldRJDO1QUGF3iNwnuAbMph49lt/96b1one6ehSsikpwl
ZqYivsx04gzVNfHORX+blXqN+UCRKz1ORlTqmgf2fIyzmtg3I1JSZyOUGYlWNMkq
G+Lsz+g0MiwSQ8Zztseus/M7Al/3haGZJfny+rObdOp/T/cf6m0FSut7wuPSFvBS
iaRzviXsy9CU8zAXRKLNiJQm1A1QUI2yuEsmMlI0wza+9TuAIn236FMdEqacqF4m
sz4lC4L/uZUDWOY5ccILMvpXh/xfyvcqFzsda4VB1NEVjLNN5rrO+tRsGmRHW14/
GC0FsBvBagE4vHOUz7v8LjXcJ9+R9bIakiuGuzFofmSBRFgANm164SIo7g8Zee9V
HsdsXO5AMGKpxBmMON4J1s5h/yOFyTvgU8lUu5zccbqLEBSMjAs3jONBMptMWaN8
RBzSfU/fvyMAI43R0NdROHkyNyYpt2DGL0OGPz/cYIKkRVLzyM4PbmZrhQES8det
lz9UOJv7vc5aWmnptXFUm3tjNqLf0bns4lap2i+UHpCHRVMaCAPO945qCwHRCNp4
PriHHLhbgU5Ym9o6XjDyeTFkphnnoQ0vwUcmiddOeWCtY66fIV8djPBG8pSF5Tf1
ogr3+5zWyln+LxbTdsVNtsqRf/JcqzD3Td2j/2FSHdwxmVAZDhmQryXtlRyPfBkd
DbGRXOZz1W3zZZEs5NMj5mb5MERlCgXZFmk9NFySu8gDPUdWcdvc+27eGXRaArnS
xKWTyX+LKQ/OHy6uWy00loNrYlOvbim4hp9NAUuZcnHd7yL1Wb5sFcaoQD8dSEZp
z5SKDwnh9CQOL+eE8HemjA60b4tDkhjZtxfwv9veSP4LCBZCf1FziuSR07xVDtaK
y2M45Mw/+QfptwQ3oyzg5Cq7igWsBA3oFMPV1zv7hFCbFYTtdHFU4uL4VvU8xFEu
oEZ0Q3ZH+et/fS130KnrbhjWzyyJ0JVFYJzc5yymxszVjRTGqK144O79Csyge6n/
CUPzxi5HfF5nl7DJ9udozwlMtvdRHvNPZjkrYUbpBds5Iw1u8afL5NQ6gtaK81Q6
z5zrTh/fGBLfGbpSFJ8dm2jxd6Vyriq41azTxtb8nbKLapyx7WlEkGJTfed7ofsi
n7dSQLkEdzBT9/KIQV7yKZ8Msk8EIcYZks+OCKShNwWUML7QfvD/55FTQc5lrxjO
DjkVcrY2ZvgA0vhmYr7L+s2ZXNymaQiz8NveI7UCZ7w1ICcMFHrDfbAKnzwJ8E/m
sDT7iwWPVHwMW8PMht6dFK7etHrHjFTc4HSIR/2K9fLzeLbwIV3A3y+Ejd3BZuMv
uw5UVwDl/r5A37GGK56bnYYpRysFR0i8BxEysr0uAsvPdnCtpjKw0cxPl3OWs8ZV
/KOrpoUR3HEpo8VL5dJMYtpUB8imkpnHYBNlpoPm1LG1R0dU7nWkG+Y8h7p1clTA
7kXHKd7EepJPx3kJacJRioDkNUol4uoaHZdffsHiyjSRchBpcAiZmrK03QSS2p6/
D1P+xfXZ/YF8oTi3/48xSJHANu21+S1SexbjA/sZV6cq0nubndQKrTdpTkHHt/jl
3EgHdnrX7J87lXAAriR82zzMgckMc3dl6ofrG7hZAYWQTBojufE/F97TIOymik+k
S/sqr7KXSYaDWemEciSnTHMvQGMW938Bhdx6Cb0pBRnYt9E77nj9DvJA1sbJPnMr
x8LgVCg6j94Du8MPFrpgpOQAO1FcoXFMBLqmguQHo7yKMaHoA9DZtNnWFdjQ3lQX
JqhgUd5ZhfdvKiBmvubgRTowwMAmrgwOXmcJyaZ0BrR/5UA+JDMkOuZgqnY5ieVY
FAkpVcp80RWxYjxki0YH76C9vrnv859/nwM3wmYYTR+VGax7jBJzesLRJjI0z6Vw
p9vMIt09BNi+4tlZ9nYimzF1zrKfMv5kUkPbakny1xTgIRG216FifHEggzaIweTR
Y6jKTO1abephM5BTTqzNiPXVoCp73tKBZT94rTMjBwnb7ZV3XcujX5ytHavYNY8m
SbmsO32B5HpbGSkmm/OHfqmgp+xVVwyByTrLvkw4xFvu+IRzDD6oZwfryWo7WIfN
M4woN6h4TKXXezm5cacd2s8OnhgE8oBuzOC0/m2rwasnWVZo57cYNzuTvTPUozSj
lM+LW/Axt9PeHA9Svg8NTowfAuBvGtcNnD6tN7M6SkMLe4AONKqicFFhIBxfaEzT
5qABggp9hgt2Vwd8e58862ylLjB8CbxmOfIDYAuZy690uzuCRAMDGsEXKpWHiZ+w
iIAlXw7pvSdMf1ZnLVT5LRQz1iLQlsQq843RUTqJlqztc0cAe6HRn5VzSif4m1l5
iNsB5Cld2IfIrkN1uWFZw5hCoSns+q4icucpjvlncDzYUJXuC+ybLej0KCLN97BM
O/yXC81gPt1TcFcHHFnNLvBwo0uXN9TPlDOCLjG52klH2aVcBZj8ijRtP/QkDTwD
5GpJ4eDowoZLaSQvOBT75iSwldIVlPznKptsCksr7fUT/g7jjdVf5NfIhGi1E7wn
Kl8G+TljPPdXHwMzRAhJE0qb0PXYodlusGRc99AHj9AYWFVNL8befdEkLSbtxn89
Q8DneF9z4wN33znjWX8PMfQ8kb47jlli1hXHqhbfK5YGXwi41t5nG37tgDV2HY6t
1j58QPMW/WAHQTOj7eR41Ogc8SVxNDc8HYvHyAJGcfopzcTa+XRBGe6CQq0CKz06
HZEg7dR6HDwn3Y/rZnp4aFRWTKAMsFKr1ojJGmV0hfz0JdMy0DzIqdF02XaezodL
2B8AQudiHQoCfOuc4QlxWOCQjKMPIuaBIEAXhDeRCEIuc1PRkRlR0BWJFY/4lgJU
LeTsi2VDlzzgE1SIhVyltgdA6OIr4f/jZoKoSvE2B6Undu40Mj50lNFvLkG8Awi5
KUTeQNwaihvnAupTgzg0MxoUFN9QF1AVOoHwH7Hltm+VYOUBVBDOPcmbaPNztqBe
VenSdWYemi2Jl+atFK3mB8Wrq3fN14ot8h9A68oHs0LYqRLivqiHYAhsGDJUM69O
BXDzUWeNr96zNdsfwEjfYr8gpustK4YBOD1wnxR6FVJQGfrTcqKXKGwUu6W+RpWO
VjiWJ0xZfELcW+0JMZUqygtpOQo2u6S62SfIFBTl4nRFN4ceWyxOY9UztR93FH6l
wqLUBwBAyA/nnexzE863xXhhhmc6K56x3j7WRiRKNl1d/x4gwF1R2lsYyUdJOuVZ
z+0PIhMTOpiOr2fM4zGRFLXdsTKS9jG0PfOMv8bqvGZi0o0AhiiGvldojyOr1A+N
rvLJpSoS+dghFM6OJMX3L94rZ7x/Wyxgzhd+xV38USJx3ww76SVKTWv+iSi2Mnd9
z++RcTHlewPEidB5KmV82gbcjfqEfdkfC6ntS2mkEAN4aFLManXOjAqYAu+LZYj1
BtdWtNyRbJRcl7JcXJsB/zTam1ECD5J6SOGSVaejiZUfLSzxn3/YuyWvVKuVowCe
6NnZf70kM1AdEut01KBFgjzKGznms3RvKn4QjZuxMe+SJDSFPSjMBQuNtr5OA7fI
AQIQOycjHNb9A7g85843jg==
`protect END_PROTECTED
