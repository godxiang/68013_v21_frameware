`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ossz1Yu/wQ6hBw3FDewRrKPkbzfKlvQRmBUGEDlKYr1V4nVstWcoTfJZslJberQq
h2YKpHEwkIdelZ2gaZ9Sc8y0G0eANkyWgLRD4g5nWrJh9c1VEPnRupRbHc+uHYuj
SKo1nVFlMZxymrl8xxXW4L9DIIpz1BlJ3pupBLIT19CeKOI2qsN6Rrdike15P96g
klLVwXHqC2i9W/JwgpgmX1Yonl3rx+O4pxgcYczssAc/cGiEHFvQBXO9BuJbCp0R
Eb4wRku9ztpYCqzzL+Hlas3KXOu/H4qM8iOlRhJ+JD7tZDxkxnnlNB952qUi7axG
zUF+KUKSV+LJYAXYpVHO6nHUPqzNnpFUd81krLwnRiWoe3bbYHhDJSfnolEf52fR
0+Wmi6tOWX+rTJxqhGc4Y4/rU5LfNLvVuQ0KL4gp4tPEnM5gZSUqhwMyBfP1LAyy
Pzh+n+EEPyvL2/6QmCugaw==
`protect END_PROTECTED
