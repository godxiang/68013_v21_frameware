`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYVfVoUecWvKVTU/B2ZZc9IELbSOTVGayYmXQgF8yQlJ2GtCccj0SzRzp30oMp1L
b/IVpUFzOGpk2ZK6V4S4iygXHe3HF4Knd7uQGAb0R+9GpHmSa3KmTMnU8Spck0VG
MT41oIYOtz3dRi1UjvA5HLF8TovWZExi1/UtemlasMJfh9T1v8/b8si3mkiJ+Inr
FcZmTqcvtn1+9sGYpIZfBaXWNe3My5XJCAe532iVU17QzqJ2FxK+IOvnPzefgkVH
0qkOxe+Rtu+jIjoze1z3CUgtWfNsquyhHHANmJ154WzVIG+PEflUyUw3XsIOrPVP
IJh1OgFc2Z7qVUpw5vMykBzs3uyvauy3oxKGTmjsaC+qyGWXV2GzF2yi1ifE8cb1
46YTfmvq6XJ4SeviDqNyPQPeIulK4NfYd3p3gWkjhmDdRQzG8HgVm+La2V9RE9RP
fAzsW/n7vkvFSD/lOjPFJWAcMZZMIp2zLwKkFkdmumDdj0Vhf414tX3sHdeWW5f/
rG7S7btbj7rzvdK0rxun9NKUnNWQT3tbDyWcXvMxN7wxBsQtUxgyNGsiCDNWfqvg
7BvboBnw+BD0Ynkg6sNAk6BeanYwEJP/ShDt3PsVK0pqQE+TW2WN4IeaBfp3CKFc
mRejE5lnPuR5gyfomxs01WnHgVXSyCDpwKxI5HRe3KoYOI53SNRZXRhO74FGVXAH
9x6E9kMMT+N3lPrSjvqtSvPuN5807DoAjB91s4Sx6IwVaIMdr8Ou/Pd0K5Sryb9m
ltOpfpQVLjbazhziymP6ORiLyZJXBp40kuxHup6AXeJzoFCZlAdJgWpJAV/l64q8
cnbA/+f/iaMRpP4OdfLdyMLBPnBWGiyveldd5F7r7dtz/RgIsOF7SMIIgLd0KluG
G2anJC2fLUOMnnMp47fs+8BGmeGfjjp1HBBwfVZ9b0PDbpR5PrycU9I9uXYmWhf+
sq1tEVukxPMpffX7aWqnJwqmHJEetuUqAU2ly/kMCvSedhmQLd4eZMWWgleHEc/Y
WoByychcDjU9T7ojGFT98vAQhBpz2akBQ8Cfo/f5IJmpTHZxKGuBvC54pMe+1U8b
1pf4vX3cvOszY3DTmywj8RvBoJsD9X40teE5VFEIKSHZGGAxtMR5SWKpxb3kidDW
x1HXknkkJV4cTrlGlj7nKT3HXw9bVpSy53ELv/uWsYlDPIkjYz4iLbUfFO6AVe+8
M5OCR2hBKPRVtK07QGjG3YnaSKFHARYbKnTldKqOKZy+haDeOn8JTox2BuFjOpCc
XhIGQLZIrDD8YKLTRchJQy1TLrxZTHHIQdki5wBcVS094+rkME/85p1/Ms4Jue8u
RtO7z16IxVObuB5vMqcskD4F6BB1pjENeBcYBhNpdnGr6EnAgHehvu6q/dk69jFy
iacaY4hoN2SbcyvB7nKmFkCwaiqObk5CTfCscCWbuYjSacDofPlXswpSfpdk0XOc
XJadTjqFGafe/Je7snpyvTQAQg9i/6TLyAuH5IkWeKH7CyUges+sGWkmEGxsVrOk
ceOGDMiBvVUob7bptgI5u4VYJPYrVQHR18wOei1oXYWR1skRvkPoTYUE0FoX6AS4
yjaR3b6bgz/pXzEeGc4cC6kn8KDifNOT37e3yP8BZf9WqvXESsntJ+YEGswXc/AS
UEdNW0CN6Z+D/PaOr3rhw+NEUtmxLdmXw3Xg4e99I26tcs0m4fgnzUWowHM5uiOb
97Er9thEfvrHkSkJ+NOH09YfGhmM8IkyrLB+d45IYFRqGBHmM1RP+5dcRldlPNSA
QMjsQmqRz1fogJu0hOVeWxXJtbD41woO79r+ep4RtEjMCBlaPs06w1nNNq3RYt/b
Ko2xGx3h8yeffdxMayrQnkK+b8M0KvVHGbxLkbFQfp0IIyWP2/k5kBlFm9HePD/g
RPCpF+Ua8SnKnLeFDmAHHZhSMFzwPa849xrnRNyWqTFJBWngJRz75YxaHne5GMB2
CeTKO1vxClxRaLpyaN9RjVjsgq9R9EvNRl7fl48cx8lRC5K/jGDMVa1NlB1PgC/x
Xl9Ue0ajkZJxe4ZUVhEdWXSX9/mFG6oulRLtE8WvmXFrURoUpcZbWlyepNLiQBtA
z8pn2jtHZwBrwne/pfioU1FzzeD9MYKtTpnTvVnRDiBXDOel/qlF89syfP6nh7E2
SX6NlsCDV3dJN6a6aq6ESr3hruMSZpnMaMgpLeO0Yl8NOVUM5uICbvAS1i/LgXTO
SqOut+DPHvveCBgNUXOAVfnzrHR4v4wDV29Q9RBqLehXTzpCFolkuGwkOJ9HBtFR
5GIMsPtci28oJCLAnOGEZ4dxeuwS+ZGY9G/08IyriOzNdVxFDIxqyP6M/4DYAA2r
yibjP5f8x8k4zy2oBZDTD71LCtjnw0+mPulzrLUfC8BUHE0kXoYNhLIK3bFSqzK0
dpNkiAfGfLlEpvgMsdgJqyojo7OrIxtkJySlrDM29iLnxbZ/aKJDsL9b26AK5q8c
92w/U9Tu+cHjs7KTyh0sFw3ippctDIPUIg/Wndv7VZAiargh7yUMUyRTZxGpwDRH
0sR09kfwLCYZvQdDNlcRpLjw6jAdvSllyQHuZSdiXxQqrRxq2MZdnmFNOsmSSrNR
qf82HXZIAhOb4X+SZAeUFlER+va2M7ELcuYeqLm0qBb0CJ7hOosVOOUbZ0Y33NXp
vWlEgdKGQVhMYaUjDuWznlta5X6kNUTVPIBJyjhuGy4g6/DJuwSri4tMPIX4PDpK
/KOm9FGha2N7dcJMd6zwAoFQv02Ol9x+Lmy0V82Z9HpGHbyN9BIuCErV2viqO9bm
s5e7bOfu3+8SD0w5atE5JLPSG2zSOYN7e7veRfIhTIfPWYw1d2Iiz6IQ6Spc+Ktr
GQYBDajBq6uDBT9MM7cseVSurFCy4NO6jrc4bJTv2GpgSWo2p21kG2cbB66eNC9L
bfwyt/qZVNppCXcpiFwLBaC2c7QMcaJsLYuQX4YUUEa1BoLEj+GJ9xJfxNiwrsYZ
SwtrmbIAXlpZHJrXvJ/1pIqjxcYyK4f55th8OnDQ4p0PLc/G7VwPNi2FD56Rf8X6
/KxCQTGvYvCq3Q0c5gVCE1PfKrhqQVSRO5r9ctt2bJKZJiiXRfpFY58angMTEVEn
/5OJcSGLuiD6pKaUloFcLsn7MwBqKX3lFlBgQ18NaBEI4y9ThNyIJtjmfpx9iAAN
wjPrAda1r140xBS3TB8aLEN1DH/O3O5lyQUwMOMgByth6fczUYs6A/AJRwmqyZEk
7Stoaaiyq0Wm0vG5Cmt8Ns3N4xtWTD18CJW1D5C3StdT1MfVRzzXBy/7gbH7BGdL
NUgfIrxdMKdRK9YrIXFGizMykzteXcEKknJ+3fcrTzQfoF3wyiBPQ+RL8eGltJ88
4h1xcQ6hvtKZ38aXYVNY1xbUBwz6WtYnVw0TmVrrwVyOqznuPCj2JZzw58xcVLDm
LZkXsa2rApoJAW3jMtjnapOVz45uXlbWYkkhq/QbGYS2aXPdXqZl/+BNKT13Mdcw
+GQbki4yBJiDXgbcw2mPyDw9T4tkolYk7e+IYNupgCTrx4pA3v+COu0xrsgPvqQ9
ePyIj6+A+C2WvHU6XMps6U0yIYPMvG6WxUeW+/gHcPfMUP/VYlAVt2qokpvU/ha6
jHK99nT/50Uhtcb5pMvQ4skCFXiVQZ+bueLiUmlCKqY=
`protect END_PROTECTED
