`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6D82tGiEJrogO/nba4hNFaMzgRULU4uOhOY69sqV9EorN9QAAxbGXSvtlm3l0ebQ
2O/UcScX/sQcoh6gGcDBRYx2BdDhmQXI5hOqmsejiQQwJKwx/f2Ds41O0c+RVOex
wPk1gIM4tfGqxB/GxFf5V1K5YtG4loDQ9XAZIl7SIDJtW5s/4PCVQS5QDAnNUjbN
VJvL7yxRARGZCtRKFXC8OyitjtG6IzZ9r8xHIfGGlrFclz3xwIAmX1wgDVuP7hHo
2BI6/qsP3g3JYawNncrFRgU9p0N1TIVcjZie7Sw2iLuEmXYo1/SoUlVCJI8tjbfV
q4AosiSvY05N25MwNuCO4PZoPoako+BziR1yvmIXiHs6YJKFyt0kD4peu31OCvAt
HpReYQsKho8O4UNprl+yNIgcfPX2NNGYq8F+Uy0gewufG8ZAkX1xUyiUG3eCwMLj
12SFAVGI/Erma0gS2QXUrFsoVzGBuN1bl2uV2uO8wnV5FuIU3mN916VsV7NKI6t4
Ej1Yc6Fabg10cOu3cckL8Qt3MxmTcEtYsjVZGtSbfUhmqSJezxWP6XYoDU2sI9yv
yypCmd2QNaPFG7bAn7EBaiVfT+AwnTdTzjteKvx32P8k5POf7QNK57lj6Y5KGLa6
zM9KaghDi8alCnr5fxcg1lOArwAf9j5Df0Ue9Uzu32WC6uUMmu6o87wOEA/9RYlf
cZArR1ik3AK6Fz4e5Lz8b13LFaaiypZXLVbHe1lRIPZMjHJ40FVvyGe2BJtxNDQ3
UfMBYTi8YUEE2I5gsUCFe1+b58p0zloNKAUDMkHHWAznCoaNmNIAzwKTK5HLvF+d
ORg9nrvq3OhVrjvyOtDPvNpJxydOb+T1YkUZCu/L2U/59lZXjFixFtp5H9NDMqH5
hzac/oGaZ9AkoiPJTi595sjjwql98GX9Ij7d8+L8g97lbjJHDIKkwtCl0/OPT08Q
wBLwcvck/fkJcFsQfThi2PyHG0Q67aEkpEc6tBi4Yc2H4KhMmZ34yGjGJ5Tmkhr+
LkHEZXobDniGEHdT2MBUTfTUw7FAzJbkKbWboJxo7tW5cdijpBNsFpWikDYVqj1U
nutUUnqst/mPt8BFkuhVtmzMWvFoA+pEjsFVl86zgF0+Z/3rW1/3Vs2YoNMa5z/L
VOZQ7o8nMgU44PQFNDONznUE++fDSxml7DaAXQHDdowX1vKESxoROEjfeGgq3ear
2vcz4HXk/iIlW9xWlwtsokaVlKPJ8ib5+Y/h5bRoRj7v74KnmUM3JPXPayl2CgkA
6jmatJ/RTIC+QpeDaJA4XigR21YZWhSUxOcvGLMt+9LP6HROzqrlgb0lmF+HWTAF
0cm+hV+IZoFsDUm29NZzkBsOfRsilh24dsUQvo/zAF6BGb1SUP95jZWHlhp1Ftfu
PUaoh+C17ve+lWbql7tD4Su0eH4mX4K6h/xAU06b4viSEqTx5RzAaVjiuOToW19u
NtzzH0iiXlXMuLFgPbbyPZPpXQzCIGCudUSKeuLdxpsgh5Jq4sdbeksa2jRmcUal
5Dfgg+GOF1a5OnyxUm0fLqOrcyhyCg5YKGKT8nw9Cbj3F1k8gnnKayxPnGaeb8PV
J8nDbYovM08ktdIDtwWQkzuorOtT0cKoY8uNCE6rVgrHJw30zKmyia1O58nbVcih
i071fRSFl7swmuNDN6kzN3uKv4OzhQWlmQvajrBxBhPvK91pX7VJilQdpKU8CfZ9
jkm5TM2eMUdjpMuKtMio+z3cAMGkrCJUcwPnLkqqrz6AcrjgIYT1+kxaQFSJfblh
x1l7Bl71tOFg3v9Hvml6ZPDncEncZvkE9SQA/zJv1zaJxwvoRJVcX4XKi/A5r8VP
b05gZ9330RM72J0RcIPqERTECf92/URoruhQ/LQ8m5lnOYVSTNBJT1oM5ggJTh0E
ZCsdUrFlY1Zi02qnq/jG29i1Ks795J+/6cWGtDDcXtLzkJkZC+U82bQKnBONt+2D
2xWAFBd22kACAvocbzUdFFoaEOLwifbfKGHQ3IHl46O0NspxZQToaDyZUUsx0nE0
O60yVlwog+sT225XSO2ncXODUpZJeOISnRA8g1Bg5CUysTG2h4/y7Ke3KtHZQ1rm
hzaTSVmDDVcaXGDz3C/2NzLBVZ1IEwvGQxdL+dqL9g10V6IfrlTGCg12Uklcnf2L
4UCLT4BskrxILnenuRhwIfEEQSDdBEUU+G+t/i7suiAIjcc+oNAijHvgudrf4okz
WoYF6HIwSsFwHqOrfb0upHOi5sgFNaWGcNdGXpoGEklE//tgirQuJtagxo7zWQBU
usls/wUWDLJh5MTv752u/ddwmufbJaQ5FZgADAOHNUyI9ieX2FTSKwwacJ6IPxdJ
syNL21wXcVxH3Zo8LLcdA/RlRq4SopRYKmXZte8dr+faT+XdkklhYNP98o1VPNMl
GRPUa+yMGCB04JPArNPE5r6ZPNuqMYSRZ1LgWcE7f4aOm0+a5H9lzmzxISUDJNKn
ZXMs8zs0JFi5siXpOeoM0cBmqMYZpKtfD3GvOX4Y7+AeHNQe9e6cFdttMDNUztrp
bNTxamXfswU6LI1I3Gk6qlsgIGC5N4FA1So1l/joEP6+3RrLTEJNdNxNHNVFTbAS
9DAYPVQ+Mr+XGPTxfZzzS+4HPamC5549s+WAx4/V4/Vf31JFEFrpSs6OBdqacFw7
/6YyxyiHqgagYwj8cVYQmydnhLwhzv7S3VobynxM79ZtUu9CH3TayqcQS+KtLOS2
+9j7HOs5qkBRZNH09HMJEWx3o8kZ67PXYEBW5GDWM4mTiGzyzoTHQTctKUlc3Xmt
yqkKcvOdX4ITwECGQdz6q7L8H9Uogp9EPLwLivVt2FBtI4EfwIatm4DDmUIaGQ9E
3ElwMgrvCsMKGviqUklaPrEXvrKDTd9TFvaOfhJxQCdbc3zCC89dmAcwAVOD7McL
O4mhSAzsOoYhfC1Ry2VyyN3KfPO+t8XfK6Tmqxu+oePufQ38YXMkfl2Il9cp3T/J
oOY7PEdsL7G47Rg4evI7tdn01FJXfY6gFt7wC9RrnzNfHW9JgJVrhUiV0pA4/QuV
6uYqFfcA8R4PX3Fxj3YtdpSeqdGaiGNFQciV2GuEA2UNMukl5jyJ1VWZPQl0H0Th
Hh0yEx8RgJL8t0f6KgLeWDJLJIDbUZXkQDGLP0fRu1fXCOPzOCd0KxShwNToNuKE
TIkrtOx11PmcU344nLgRjHBvUjv1uX6HhvxqcDCMrfHsms7QhxHVFDY+QBuMfpxl
EO2GlBxOixCwTyd1BbrPEvWmm7KQAkSgtNZ4twLUs+yMgzPf0X8lV5qw+cx4IQ6o
YalXBEH7W6jgnolKVGxOgwkeMUB/4BHYy8cmPp2w8CBP0+8fJapU5zvTSH0Nbr/4
6qHDCqlXnLlpvGnczLqMZewycmUnJBYKRsg6rPtV5yt2gTouFbfdWioSNe10UTAh
pUBEeStzDHnSLta34dogX5EI63ov9SsMtZ4BIvrorlPpc06hIXlX6DPTlH/UeQyZ
UTC2Qa76q4TqM807JrmyrTraZS9yJYd+YwnX29MgoiOOKXmxzDAKv3CwQS6LtCkp
6f7Cm9XHhXcr4cFMZrX9TDGJbAnQfUg0btACbBM8NeLdlckWMenF9RUuo8Y8qUqy
xkjfl7mBDOcSp/mmVdTcN6pbd3m3xolzJrh7c+Vy/6u2YSVlTQUTUFFWl7NPmRgW
`protect END_PROTECTED
