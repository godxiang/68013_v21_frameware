`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zl+ndG5FT2dW6OHeuxU7yNoby6V67bwNklBKjCK7MKCMrr2BnVr2cElUhChVx7G6
XItyx4CHrvjaKFjqnwLrQDbKnPg6Cjhv8noDObPXfQ+4d7D0ULPPOitu41rGXjQz
uogGHglbL0CsvquQymDkAIQHmabHblfA/bhEu4DHw9IlvegWFG5m3c8QlWul+fzy
gZXElLMCuSAGzVg9zOErPyKhgAkkL887R/Nt0jFC97SfphvC7UAp+0ymz0MAtgFe
EADNP9ttcY9esdG0TBbQWJqysKSBB9O0Z7EFTINusoBRqTxAGXw+txu967mZ/TWU
fQ5RyssP1FsKhVTkon0D3ct6DvHTznARqemoON7UBVIGg5C5R0X5LaMzY7IwkioP
lq5YsFjYgIUpb0WW8pdH8foA/mMlBWnx1/wmlE6J50bA71ZfRHx/+CAJE9q4j9ty
66pwPvYtt3Ct67cT/Cx7pJrOinsfj8i/Ip/Rl4vkcwbB1VcRzIKOBDPDTIEJHzmy
28UOW21o0GYHofn+UGAU8CrJeQguSleceV2c2lexXijgIjVQS4034fTQUbz66VG/
BFE8D4iAq46PeUDUz5G0P0z/3mz7EOsxnbWNm+ANqUb1P8SkdhMuI6g1LeQ5055x
FTxoevWmdJvXMYu4xj57E0IXGJdTJc4Ig22tASj/NX/0OCmTPoua2Eio/FtL9Yv0
KTd+c+fAGGNWLgh/KAgdRmpdbTn88v/x2cvHES8OUWWdCDlH43qJzHZYg+kUFqqO
tfKrqXalSCrroefns0FOwLxyjmBDfL1t4n96+eVMf9po+JvuuYPHrbtpk9peCjnC
ECjZ8bmGQFqn6EzMjsxN8GDMvpbNqHD/5K3KaUWj9LQpxLJVn9awuDwOOYdCbYwq
2tf1eg4wd7lCOTwCRSaSE9g0HsMziS+8bR9bDNXAR+RW4X2NCuF6Q5DbD+nl19k2
ZLzeHhxw8dkIM5pwtbceZn6BXs7SDcwKyyVy76qaxmzWg957Jh06sOxAwiAvtxgF
xTOPXFUDZNEilP38T0bT7D3vjj7FW/hjyzbSmkgLXl0OnJKYydztiHUx0dkzvUGr
l12Ggje998oTJJVXRgzO9k1i2CCvJFKsd4P+79o6TdJRBzTapEvCTIZC2k+vHfNU
BXTg9MRGLYv15gSQzqY1ovXlL67v99KJtdEA+lCfF+/aNPNBsmdFxTXP8jsrT7Sv
9Hgc3JNPvkifuWI8b3d7d2KPodha7kLVEJUaDEx82raS9yTe9p+sRx1Y+TrlUMUI
okONcH3j7bIt0S6TVBETa724Dp33R2a27Kawi9AZqBxZG8URC60lpRJBWajceqBv
nlb12B8dSvg7yjgwzvz0a6l73fh8qSOPtTMtLRw/tuE/NxfXlTthUbX4ikevu0BA
R/Q49v3mfBWJHmg9gTxH8yLxmLErpU3uQ+smO/qb75cnE8QEGDbXkd4DKBkFAxOr
+1ElHNiO8aePlu+8eu2Ix/oFkwJJ/mMN+cWn0zfXLBsckcFVpGVix8/sf/VHaPYN
ylbkYlbrp5TJbv5vzm+RNL112fk9byKVlcTFVNgdjl6iR8H/cec2KsoEsdWVElvl
5IA4QyJv4FCzpFT73qpFNDS2nZBv8Cg6lOMdL8pal4Ph7ABbSk4qZxT28ZY2i5WC
Ys+8wrOnZsA6dERABsaHcsyQU//JlfxQOWXnLWJMDTxIAMrLAyaCLnI/yAbiPok5
Hn7/5QsI44vFwjOapACXGbsRmVv+0udeoP/AByFCds/vizUxjPDxLkFJQtKrOH8z
YNmcFHJ56u71HmgUyxpvTc5oSXHIe20OKat7UmTkGG1C/+lcybQACXKnE5C8mvBj
d0ONN0t76bJhGDkY88r9+cuTNdIay2crjtfbUdxLxtsbQSXRkIPiwrhBmfXHU5io
+O/EA+8iK0rR0lkmutUGyjvQeoTm5l23wSqCNlKhIcR0YcgebqOqAEw2BuLNd5kR
kxrSKvDkXhInfxDYIZY2NrveSr+j7JwpWO0SHJMVOWjWyXg7/o6xC8B+v5yJVtfU
Zde7yNJW3nwpvgtCv4Uo6/MIl3IDN7iM0pmeDEo1sjMmhrbqJ/ScLfsMkLsrHSB0
zLSY5QKy4U9MZYRUKL2dQjoDJq1g8+TvBaRgFI/7gVC0PYcdYPyAKi73GIJZUfpv
ZhGxVNGgPHqzoJ1JDwYPOUiGnFSDemqYOfK4Av65cDKhFgtn9ZsSV+nq+Ihdj9Q0
dbhElA256fZwq6GiUVYIPN/PPr06CmlxmtlBJ2w4S7tcVJjB3pqqLMiVT0ORFfv6
zlZ4DKeES7gBCLDT31iUbrtiuHWa/yLlvHiO2+I9talqMtgGUo1+sPA+5JZASic9
5E85O1524ppRIQSorWJnEDvtbAlCJnMLYm/oWM230VQab8TyJIuQqxq2iEQqSrVA
KWRqp5WOg3aU+Hs5+6gxY/AwneT6NsUvfZqmNAzShMvmfNIOkU/cbgI+YshgWRg7
A7yK80YBjUBSl+NysSlt/M5BWWCxYMGB8ltKUduijYdzKCbYkJn+OYmtjU8ipGkR
EMlUw+i9cOeVVoOQpSX6nHgTnSYHoCLcyvVcqSfKhJON4m5hP8ctH+BMgc2jCD0b
uNMTjMIBYlrEw+2j34YvZAqENcTuc8Dfod9qPXWmPZ194BMy0RhDKtYPHKY7kyxE
LrMn9J/vE64G1xGAZsh9KM1BrDWD+l6/mdzA9nzfNejR9ZtYS9QUvM0jdhglaAJ7
Ft9dI06yDy/jSoila/7oSsPDXI2ZZIYINBUCuB5dVEJAQOChi3fkwPtQdYaSq6QR
WqdItKZIUMUi3UkUvq7nw0slxNic3UhU2lJXTcjDDtkhN2RGwk3HbRONDiGkhod8
P+Mffve26BLUQg0rnSoZUYAWQt8adS69NpzgdVxxdRF5FvnuJZdEQyjjHvMsj3x8
5led2KjozxyXSxGy70JQms7pspmTsOjfTh1FZurpsl+efSuRwfoCB5mQI1Gc2D0I
OCBDJQjLWVw8rkBG5Wyv9RyosKNNHs9XXM0pUHH8EpkuFjQj5BdPW2Itm9+mUMNo
5KiDOZEDLi9idxRZ5V9SpyD0Hh7/RB2xKyZZFAf6SoYO0SEbJzyklCJ8PTYIs5EI
xnmIz3y88kIi8Zk4k1AihxdOVjdy4XUOj6IrSXRwh2UWwOuTthJT+c47Vf753x74
6i7JrOEa2JVBqBmPgJe/qXpW0aLY+9HrIlfmahdLrPl06Hkmc0AHtICQoNnnd1vM
TaPdviKv/fHB/5MTBWeaOsVAfAww+vw3dOglDyfoInWLy7Dyog9QSgUstJgpyceK
Tw556wwUI2SxvKWgtZAdIKDjISbp3MCmLxB4ja3Ssxl/HYk/tFxm9UmvnwYkRKtG
ZdwWwHK9GtuSOYUAZnvStd8Grh05cTRiMnyk8PnWETxo+iqNYUQaDURa6hudsDzq
nNs9av500LhN0xg5eTdafVt533b9httwyd9NQ34VDQpKPuw2A6nxwvxL+FTWCwRI
+rTebQx0wGZP+nJ5fjffUaV0xc/EJxmjQMXEPg9MhMvN1/BjM1Ao96H/mRFDPMNW
SBIs/XnaSvaqSP1chCrzOUN6ORhfYJYMrzNQfKob/neWZ1vWdtrqxaQNmU/E0Hw5
fInkMuATz4qGLtzHLZMQh9XTdGcGP85dbYLn+EX1D8zriAB+saatwAFK2yD0P8xW
b/6mcz7UnvrCqb7jIG22Uc29nLKc0XWYT+01bzNQURm9LY614o6Ql/zquytmkQUD
t2n1ThCWow+cvSGyDRlCiHjLy3tZs6SvxGCJKCMNVeJGGBBbFH6Nhy4e55E4Dgh4
tD+2cUhvj4MNbZpL5bhRX3AxGg+Uqw/i29gZLGh2RFSUEGpRS8IEiUNj/MLUHeyH
WKivSTlI0anuo1Kbt59895BgHMGr58x/hH//G4VnkOomTTQAw01AcSDARkAe9OX/
TluHNS6MqGt4hjoiIoncnSnNWayKDAETPuMmRSmnf7p9TxoTdwtqevtcPrq+4w1T
gYQ8RdoR0xGQeB8p310RgXTehC9deZ9hE3vY2T8dTtWcQemPdLMAgbNakJWltcTi
L0GlhoGijHJxT01yYW0R292wSgg87zQqQqiw/GYFiWg5HN05zfg/cY+4QnNEtXvv
VguyP2FaRtcxuVkL8EdlguZgNJ6NQvHmX2g2BFzPL5id3s0WW86Tax6+Be21aewb
7FyekrwddB+MsOfdsT/qDA/uVxsXWQjKEZz0o+ILCIQF4uMswkhFHRzzidPWMeFM
ZFPJ3dFAfqWhRLzfakJYTfogWDFwcgpOjjVOW6zlDtTOtexFLCKH8Vd9hUqYiNz0
VirUw6d4cT/TC4W90L6o17aQqjvvbMiApFSLLsSXmaLTm6JZAzo6kYcLUkzn0JmE
8bpCWkQEgaVwNtUqdlQs23OWB6x63O/k1r4ymkhw43rYR1yCHVDv99vnN/EzyqDC
Vog3hqMN3GdbH2uUrHU1LqOdMx1ESbbm2auJrykI4gG1AdW8r0sw92LMfjCGUcM6
QWlMtCHW4sPMkuLB9gDdWYo/IAEiNQ4z9gky1wyl+r1koWjwt+SdKrXPoVU51ZJH
2kOy95ZNakEHjo+fNuGdwHhphAm8awK8I5XaWT6RJzmbNh9/cRoD5B13CP/KBPz6
DAC/yxd+4J2+EpAkcXZeboluEJHMGwl/6Si51GBF3YJYP089t23tp4n0RPQWAuRf
ukQe9o+d8i5UeqNP546Ie6pV86DYroMjTgjHVu8ynjt3Fff9BThOewVtAcee4N0y
UFqLP7NaQKTXwcl4OrRIItgeb8/h6FHODnF78/HyFuD/5hkfTYSCk2h8L86L8BfQ
C60KaEzZoOKmQB7qmj/hfhylJTWJRm65FhS2JUmdYCeq7GNp0k1EtDEq2nOhLvZu
sklEiJOXAHttzp45xRdp/A430Lnf/+/iKp6zPgjN1UMkDrOZi0vdOwRZH5hB1k6y
9A+cI1m6ptZU+y7J2JK/mR2nX+NbNOX2EMGKZu6pie8B+f04HiAkSvzqaR8fvqVq
12MUkTbrztCK2xsI6Z4UaevXNGhJ9GJsmRsbJhmot/8R50voat4yoBcFNdWubSix
wpnqbTsm3XPf/Uqq4qgJkdi7kI8yc/zdp9Cz6xTglmMmjtmHvN7JUcgrTUYnBz09
8Pm9nJSjshhFX0S8sy5WIDqdZYIwTswxI7dCXtvUMktHRglu+Eliw/yEPD4q57/5
SaeY0XMQlYSk4+qg++gcEoSyrqCOJtOToC0FWM7cJsdAcnPXINqUgf0vjHBjZ6pG
1gR5OD9Vb9b/nfcJkSpDai3Bw//D2RBLNCiAPqMCd40fHm3ufAeLwtDeTeP9qr3C
TFZIeQnhiRQcp3LmBpEPYewbzZ/pVBIVi1myuPAbUvTqnDOQ4TuyegGy4Qpj/FKq
oB9xygrkigM2NkNOt4x8brmLJkqFCqKESYB2T2jVySGYFK/ak5jYuDCXTyRuY2aq
nmsltwsqDDdTqOgqJeqqy7Qoi0LpsHR3Amu5KDfHd9v7paUcx5/UqI1dWLwH9vVv
fXqXyL6T78/Wgem4KY5PhN9hf/5a2pVDFeVjf0muJljDVPpd2V5sow2PStVz5BKe
9Mz04ELdVpm754VSguYP4aEanvv4YC6GhO4z2lRAIBZS403TN+D5/RM5ljJiCMZM
fFjSrFTyZX/IhdLa2vxhqk4Zo1yBBu60rnQlzL82jVGHiB9gn/Z+AmY6LXPJkvKC
eqEehAHtfqcdB2R5ZCULcdart6a8cys2/rykHPUFpmLsp/ZLAZAq0icAvuWLbGiy
q9cyFeC/6H/iECZq3KnulV6MnyrG4wVTRBtcjQ+Emb5drAP2Xp4jcc3lKYRwbten
BYhbegwIIetVZ+CjkidhGWF3uyxYRC43JmHcxu+/45kcljGAHAtS2+o3Nj+M2WdQ
ikLRzABCSvOBDwDjizubuYbKzIFj4DNHWfARAOuuUcZI173bUB8BeOxlL4KPMgsg
94PH+MbiLFK5ybWoisOG4Eg1msHQcBzSBIUyLex6M/bqYdazrtFqIKw4mqJi/Y+7
CrlgTFRcUnPPWNedcCD7oXLQQnTy9pDh61rqEU/b1R3MX5UjJF1RM31beBsUh60R
MN6arUTLid6wh9Ll6MRBxjm1CTaSCu6ugDO5cUA7X2FjB6m0O833rmGlIwkkSt0s
Mo0r0dxxQzgcU2osvOuLDgjk3FzLVCNEBCn+gub/XYU85E45gLIBkYlH3Ii6jCPX
zrge2x2CHhBunupJKMUrNKvxc6VeUSM3lHxsLUWNdVa4zpY6EFPn19qZMCTVSQPP
AUJ7tM+LgOBwCGbVHTD1l08ZYh3G4I63i3EO7Plgbj9z6Rh9fAOW+xrcPt7RODPH
vGu2JD8Q8jlrKpAdpW6X0X87tpo7VgVmPC5GEeVK9TOPcZOR9TMogrFZBt+G0+JK
yX66hYfAqEUjYcX7WBviFc3Ym4x+X2caKtWejon56bdZ9QL9BMek64DguPfzt7b3
RXILIskVVczzk/HEpyuBmdaSk3eJuwUSw5FnVb9AKehA18OjiOdd3rFi8BYcNkRk
wJR5DeOxrQKl+q3fALJxooDu7ow7K2OXNQxCW1je+lnRvVeLWmv2EiAiZ30cDwFI
vmo0msZX92D1SnKDgXbM6f1w5oekKj0vd+HPmgWq+/HT7Ec+9+2SW2UyLGndABDj
pgOC12yuvej3XFLIYG7sJB8NFNueNfZK1AoErJPeYUtfbTQGaJP0/MR/RwLjJPbz
C5EQHwYwCENmhPNphy2bphLb1U9cYJfRl5lctEwOIy4L62WIpftAq01sCcBoRceC
VQ39TchSv3GMtO/m5Mm23UmGnip3xQ2lAMtVIRj0NKvvdfNAtnhG3APG/abDLOUM
GwMa7809u3SDMopPxGLQghZh05stnwdVMv0lDsws8A4IHcbd/NKVvBtCGCWNP/5T
At0az4OBYFNJtU5AG88Kpm4Yd4baw9TJIJ4YfSoA7cT6br22yB0QOAHao1j3nD8t
ahFegNBp8uSKMZ6qlxXCl7f6tVgvy60pzJYjL2kK7LKh1+yB0BUxZxb4Fyf4yXoD
kUAir1o+e1LAWRje0ixOiBnen31apDVFgMyP5YZBxgZZtX2AFNtknOqXcS51YrvA
zIBXZCkMni2j92aGHTIVdCgD6al7ZsBnPrbUcEbkPklbpGniR0T1skg6WtUM78je
XnZZ8EwkXXNc4qPwBPNXfBsjwIgNwEAa31gh5pn5jTnUNuUXvUE8xzNja6fvSw00
P+e8o0Tjsuz6krKvd3RpEcpohlWIUVL/uv+N45Bgho5/ysSk6HZnPcviNRF7NjWs
qKVz8IJ7pek2GNVLxuVysXf5DD51QbSutslDT9gcOavRamm9P7aHIXrgaH6VICIp
8uyZRciSARk72Xye7kiYGlMqUU35WGYQ0qsWOJwC938rcvkIoJzvsi7+ijkKCjss
49EaOcbyUdtEgKz9mRmclV9PTR9nfX3OJv5/OS44xv3ZbcfUGojgo67bzaySLFhK
400+gdlGYQgaVUSCCyU3ltATuiVrk2c7WYj3/PxG+tHRqwbrP0DCy2klEGcQSqX6
K32bqDB+bfas6QzrZQgGnK0uSufLvkuX0iFIudMaWm7dzzRmsiqQne4qPsfdiNvG
e0to3N1DcdgdEZUyVZpEKgdwperks3/5o+QXNkb0uyQSjtvpRQHJLuT/lGyNKOu2
95HCv85clXbdPvL8R0a2l+0mPxfpXMormvRbP+u+mgHLAqHAhZWE5JBXzl6pchjI
/udfpSEkpytVIzrWaRdjfTt8LZGZqD+QgF2WedLVtvDubAehdG8zn9ndzN1EFOQJ
OEZBw6/lxiMYQSnjvb2NEscaEEnIML/W3dp3MzOiEmhFWGdHYaUUDfqPwsP1YV+Z
1L9UjIgbEAgZhN2kG+ffgz3ogCwrfi7mk3yyKdcvGy8zZfkUAM0jJF0qBkPFrS7u
M9Gs0ZYWzkFFgjbWbVQtw1rGegKKitGVmiUBybyCFztIjdHYbs+HGkU8+5TjEuDU
v60R9jMnI+91uKi7IcvJv0bAfq/Pcx0cC3y4R/N+1PYPqszuLCCU2aGdaEbLC2sl
r/RlUVpIcekaObViiZ0vNaRgAFO/hCxxllet7/2PwJ5sXAKLrHuVJchgLpmzjT1g
9UPCUMmT8lOpTc1Q8WQh3tlqD/dDSjMTffuHSW0tppmLrmyZqZ/t8RFyCUFLoGWM
rTxl2VGieOja+2dRm3zUWSUmp933Nhp/6wVAOx2lOGaFGzkSr97fx9rsr+lXuOxI
t+F2iaaHL3kZ4YCOjYTxXUPdv1RsZXfU6p5Y+e6pvTg9LY5o3IypgWNmfsoJs7PS
/rlzuf84qtFaVFwaosnHAKq73SninEw0mv22c0JJ9Ab9n2v1LB4iBkOzhyW1YN8X
Xtzr4hwbVkRqSjWLy3Y1GMR7u8+ds9YiV0OFpoD7WMz6/u3NuN0Z4UV5D/G9+riy
yzE6hVCyVqjgeNJ8XeNefeVsbDMpUz1lUbCIflNa4RN34jpz8K5tOucBca7eZ5UW
Lb1EjeeLqWhe1l5miQKWIwmM3pNPOYdb2Lfl2DIK7jXSwWkEQfso/UVPFqKR8X15
bSTklPDkwxw/z7PSNqVIAvS8KBJ3SkysyT4QPtMEkfe9581ln+mQRK1QBo5dQYhx
Lb01FwXsGL9oBozTvPEHKWqByc4fcMW9phEjVEexkjCjd0RdlJGlniTlsdoyq8tv
JMitvgus9SCoTLJnXuH1bJQxuvbNkv2DUr0NEHja5xqxSdhzNUsqLZHXRdI7wp55
kWlpcej+tQ65HaK3mn5fkEJQ8tq+cMq8xJIK3xFLZ/8j912/u6q5M4EoPBo0626C
8+jFmymnoTuz0TQ7ZpuDUt7hVCtjqfG6LMtxrqEERhbZ5rskLdns6DruxM2Tv78s
RiL0AVzkkx5nQtnnOJl5W4WUnXOMJVm62HtbQIOnak/TwRSjjTu40vyMrE/0UbFv
F1L9qzhhY1qvtO9jmcy+RmJIEY+dOErtnXmNXYHr+FljoPVOHOPs84bamRA8FhsA
HZyMBBCcAQyaVIivgLzSbSt5Lp4vPd8Mi2Etq3h4gVjygdKdD3SNsQzuWiunUXAg
lsIJetmI9coY+HLr672sKU8436hNIBDIKVvPbGllgzI7lNNKz9bVpZng/T0pvXhd
CPRMDkcEy+07SB7GO71OC3hS602jnmXMTnZvH6fqv5cSh/PXA3sk+RDoYbppF7GZ
3qmpMOp3WsauMJIKRQCkck8GcdztSbRpwN/GmeHegMwm8Cov9sVu9pDvD4/u9fut
+vUGM01abAhszB9bTqIXc4i4yUT3zk3M7L/L+R2kqlhg0HBIvl3dGzyJTubtzwqC
tuEpKHqTmvTy1tLhmZZiT49DuQSA1yW/iv2MVdv4TF7sI1FnY7Y2maY9K2qft39V
9eWwgrfqByQoQfELslZgzUHOUsQM/7laFyXUtGpum7wuCKwddgJEb1YtSMPu+fLI
ej83zfYCu+iauGID2WpJ4fBiHeF9CYyhX0pzLqMszhxA1Y5ncK87WSqWPvLV6jlW
HAYg1d48htt1dzlhiOTLC8Yaf9xOZZH7CBfdEEqScvORXYaucKQqAXuKUwZO3C0c
Hx6XR5UKaRkSYBQKt/sInyXXsb1iqpbLLkDl4SQChAAiu0zYHnaXH1Phf5NRvpr6
9C8Mj0A7QnXlQC0lenyBJ5dJv+/QPc0noA0byqLi8fX9DdNp3TllPz54/9y+pGOZ
laYdJFOPSE5CJOzGXcMKDfLbND3VNI4hH7j4U12V47CHrvX9lAowDy/no1OZqFab
A8yiNY91hVMDHe3HasElr/7b/g49GW3KZK/aIA9bRjIMGu+Hvztkxrkrpxgq6FOO
9/TXxjnpKroWTLAd35ea2efcoIsMtTaTrRUT0sc3NQsv6FU9PaY3Qspj4tKqbzJA
+CRw6NQMrI50BQHo3GQ6sDBtPC3+rnLFuCEICcFlJKEZAE/A86/VYDn2hQLyR2dG
LAm0T4tEyvWzJO7a5m7l3X0XekDFB2UlPRXDpII20gzl5dFopXIgxVJLHVG+dOsN
jHwVq/+QRLdIHYLWanFaAyO2xyB5K+6MoLOdvgPcqSdzVnKwZEsPQqvCLK2xnWSi
bRlekVlyb6IRDv9i/+wLE4MMwkozUOyMUjTc4ZGxjXZ6HkNnAXyuovo0N6Vehw/O
Kh6N4HXQK/W+mUX5u8abBJjnNaycr2I9K23/rhAnyZ5BvxRuo/+efZMKT5bujE/B
9PlWd4tkh0aPslQAVqPihuMbZKqO4wAvajigo/I3niDSpCZS9nmPUIPavcvJzX5L
m6nFeTvxUicWzcTcJSud7xWTUTlfUL+cAB8OJe8daz5HqTHS0znf7m2CbGJqbtl3
gjAfSGEYjJn3d/gY2L4pxLdRxVtYvt4i/z+8YCYSH0Yo0t6AfkqumaRUyHoDkgzq
9rnrSht6gQEvfFuOmsURTUzoAqY1w/gsjKrAGI886z88r8TVAdoGzsHi0elLUOml
qjnDY8OIed8gGI/Dv+Q+URXi0p0eX+k2/PaveePqaiO3y6M9DZuwbK6VSccq17HA
pt66Krqf6dafqMcFhqTqr6yIhYkjYDQd8CMvNsbVarWh399kDK/di2g+PfDeq0wf
hE2xRzdluAL7rjIehHdDOSM6rJSysUBE9xbXyz3/4kj5Umah33yU9YjvQE4parCn
J5PR4bbgyvRG7GnBrHlFHm3CFQJMVvO0uaR2s3ECOX0lk3xvl0A3YiQ+iZeo6PkB
G5ZRotLXR/pmbkFl9qDhE/kN3xzX309ZHvH5y011HMFaYYc/zc26CoDbD0fwHckk
yQiE3FSBYKd2zOvgApURFQuPg23UYPebOHYcg61tje6J40z1GTlWGWQJMd7+0BSL
kt7b6cSaCb0Y3OrzyA7Tw0TvtaHzROnftDhnO2EJwwIcTOA4FiwEo4Dqv+VbA2A8
6Fc0S5ll9Cs5nV+c6OVPSqf9AHU8VdFbtm5nAN4JjUSIiWikkZ1G9j6j80Ffz8vG
s0QhbzH9Yckrpu0IU/oRVudjH0Goi1ae3zDgWkui60Hz8qMgahDU7j57PM0O0P54
pwHCIT9WumbVQ78MRhNyOUy9A5533S3/srzq4qC5u93noibEMuHU5q7w0H9lXvl/
AfV2KWZsdJ0ZWkydn+MYuHQHIEnjGTP523tMY+S8MjnU5h204tmj+RF7Dt7mE/qQ
QDnkK6NrUOCF/++B7cLS9sr/BqaeboXBqzPf+f4mlog/hX7M5OKv2dWUDkDTBhjj
iuv0rOd0wobuK3TY8y7eamtM5FIHPp6JHuacNozuDQ3saBPOU/o9CwPEVJ8oWr0M
J4LYavVYGD7ztP1HNDZh+2I6ZUcAAcIg87jxhU+K2jC0c2Wl6jOTG3XjpFoYN6od
IfY5/bEDoZ3ck9H9QbKbSH6szJuUUUKAB82ZisHaRWsrTHsd2+ITkEee/SVReweS
qALSXndXKWZROn2gF/X1T0qbxiHPBp4PNJRP0mVS0+4NwDXy6IEjYhFGIbFL1xba
EC9SgO1ZQEGqD8rhCDx3faNK7C0n1cx5aJMaDda/SMGjO2jNQJi12GgK/Gmv2oE2
5/gRRtLxEeZUio9UaB462mZG/sA47a60PnNwyzNpvPkpYE5Zf/ViTFXsNgR8nP3d
IxH9wlxIjfAuWIgM/iOsYmwoT2Ik22/mrlwSCvquSCS66wKgwEJiLTGpiK7vv/Mi
a99Z31JnOYIqiVyFWmtL2s4lhabE99MAt/GUhfEjY0DmfFcHfonYIM03TB3sYBu+
AxnzPh/CkIuIpIORK3q93o3QoiyDNRqfCgwACbGKhnN4bIiTFFRuDyrmK8UiClsv
qJ40NuRAymXQ34+6+flTV1SgFSR+G7ZpYEzuq7S78zV7bTP8G2y+sNj0mVvveuwg
GgP8wHG1qe3120o+IHznRLGoLDHqu/Gtm4v5IJpgqa9E2uxBkTYKt10Vgkb0rJX1
HyFaK3O9cadJkO6jrfL3ukZV6rxBVYlz391Ub2QddGSFAJ1jQPMaxByABnxm3HwK
CcmW3hQ0bI7nOyqmOeC4bs8GreweVv8w8d9jaJxAaq9JtWXAkcOXKauvVwSsyGlx
YkyEV+r0tfF9tEjo9+4+SeqOSc2YnAOBwxpuLu1QoZ2JqHbAwq0TANQPwzF2v8CW
3QHGTKwdxmt3/1RbWtW3ICwvM0Rt33I1t61SE9mEvUaLOn0JhEGdKQ75KQIaUz1k
2nhPN2QklmWdJavF2RhcH0jQkfm1fJ8Pzx4iNAn2ES+ZWh9WRPxvIyUMdymwuwHl
07bAzRZdCEs8Pq9XLl3NCvOsD7zdzQ9GoHmcAwPQOwNpLS3v5JBvjTP2CZ3J7CWs
iQ8YlbyHKMeqVYi4o1PcV3dTPy2unSis0PIjFrXu+k8SPd1rCKpYCpHC1adKo4ja
9jdWccE8oOMx4cr2vCJi/MGTC212o3QMdJDqO4Tq8qw=
`protect END_PROTECTED
