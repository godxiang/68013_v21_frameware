`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNvL5o+t4dGlc8kdcQ6pCZu0yOuac5goPWVtW82VPeVQocOgKGDauEHdxosySBXH
A1eODpRbH8A+xc9M0eztjCYwA5ZtcEPQ0bhB/Kbx2i6RMgZWazzulAInHxq3y0h4
oP14dGdP2fvHGjETiqpQjKhgNJK5/W9a1O+BC69j3wOKY2hn7kAZuDLguiV7KD3A
+g1lBW/04GTg0KD7G/tAX5wLWuoUirjGqEFwq/zQl7NOPjqlvIeN6T9uWyPuSOK8
/vFqGsQrfbtPIP4YkXbj5eOpym+JELfPNDZiV/I8yqXU0mIrPUu6i54eQsc0mnGR
yKkx6FojgHK7KUl8WxGmEr79mM94U6ud/kYa/xTTEkkq4XCSFTnVYNKqp2y74bQZ
kxED47ACRBIZxFYbz1JuYLv7mUi65EEkpFMclvBQvrJtoV9WeCIOHIkRVgofkG1K
VDQg4IlzmqGobBo0NgE32r3rg3TXrg57V0J91qYK7K97Vq8+PTAk3bJBglDd+V52
Bpuay9Rc7KNw01nSC58E1Jb2GVkKz+IvUsCnS8Ig2QV9eXEkV08omr1QlUoWWk9k
tEU7CFuT1GFHs+5KfkytIQ1dN624Vj1OUjnKKOCqIL+xaQDie49IBJcQR/IrotQA
Q+GM+9aMB3Sxi1xRIoHp7ZDXbWCRZDq0QirNZ/9whEEtnnscRcdSSrtY5mhkI6GS
gUe0Iwc8saGMGbYHnMVNsDRSFsfZCJGyUlilKmW0ZP/EJpFl1+78oB2X0sqvtVO0
8V3PsaE595CRHxBYUqv4ubQrMLiS4brW+33xPYs7yYJ9w/cqiZf8nIoD/QSML7LN
Z+9YwDE6+D9ASU2udI2C7fq68InwQv5Xly8FfpqTUnwjJOIj9NtG2hfbsJw9fDeq
rQTlkPvSycDuhjSVzfr+7tYNHtpNTD6m+o+9b3wntzc/l3LjT/Dc3sBlMF9bMXGy
4PC/057WXXr5lno8xzrDxmoF+owtxGalhXVucZ40YM+2/QOo4nX1QQQSVtCbTCAl
gTdkLy8CoKL+yRbI5nXHPF4fn+JLPweun+9s7kpeg6FL5WwBnoRB65hUfwEHZ4Nd
21JT0B8eSBpLAi5DvDAG96CYGanuoWwr6vu0g6Y1bNY4I8QkpYtSbkKYzyzhW+zq
DLoovFvW83kA2zdw/gWnJTaHqwjXWrSH6c+tuX7DYJTau1vFGUVG1YPUlbE6kjmw
Sx803jWsXdAsF5NztYkkZr11j+MkOGl5T+Volum3WBLXqUh1dzihV0x5u/Izfu85
CA6FCo6roUCBIlzoRcPFE3pMV5uaB9idCgvQn+1OeA5nQlg6K6A/FGqVmCigTBkv
ofVyUMgDKUm/lQnSQXgkdWnU0awPgxkMbpEJsJ1zVUOp5SKC0IeQVpHieCjVwM3h
ZKh1Gj3TAPYwq2CWjRiVgIJPCUPI4b6Zbi84Hl9IwSvCt+S4ymt2lXZqIDDZ4qC+
`protect END_PROTECTED
