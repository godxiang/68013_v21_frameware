`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAcWtmq3caW5SpNvAad+YANzYvNr//Kp7VBLz79RbOZlSGobJzPnKIYTGfJZUY5Q
5H3y7QYkAyau52jnAbquDN34TGaSMrhhAjL+bspu1Poh5eNI7xiE+jPGs7LAxMmb
otDAv5wUN+8L1To1GpqHga14sLoqPWNT1CPqHDMsu6KMHVBeQ2MgROGzvgfxklk4
2Z17W1SHZai15jDwD0CVDPTbAmTYlEinX0IWEGwqiKuPvWRueTOjMo6Wzc8Phd0U
dbzqXncjiZZMmxC5qqdYpy0OKDFawtwR/2tC6EJx7ukgaQPY/UreMli/LOcnQ37A
4fF6gjUFNsbZx1LY9BbYtour/qY61ngiEIX8S1OWggdMV8wHiqLjCRgzncaOzeMP
/WNepxsJmf8NXwizXBjHf3/vFhTpCYtgmb2VWNf63mXD0kUU0qDzveIl7TsOZRYG
EviQJ/nokrHOpFarp9NzLw8FWVZwUKinfC4o3j8HoeGhgWi/Vuk7CH2cK8mX+1NY
keuMu2eKQ8YeusE2mjdQzDt4LGnzkwWOMPoVPP4F0h8+rFAPipkbsOCDn5iOyRhz
CFwNqnJLYVcIeqCjMUfuW+OgK6f1GE1rk2reGB+lesVdx8/3dXrS7+sFz9EizGTF
WMnkiRPY4ery4bCgMUlYnib/arCs0Z+2jH94250ZGJhi/RMjekCHcB4p7bs6+/EK
Y3nsnqSDQoS5sllhtmaiK401k8S/KN+eBcZJGcaMo6BzMNwEX+WC4qM3krVNgyBD
Mog7YJe1aTr2LGygSUI3DYIz4HhlgPArxaKcvLafuJzonY+ou5uti4ZLlndzucIA
pcH6OJaIxRVODHbmmbzBp9zaX0zeX5r0oIK9/Hf9Q4xPj5I6ili4tUSCKFn1uIcH
NlVxSFpwPtQdClNejvpDTMhQmH0UOFSMiUexMoeWsSF+X0DzXGQfSUKKPN/5iNoW
7fR75qCKhK8+DZPtDAzeWb8GbLBLIBtjcOUADhrbDRVX8Bxd6BAmz+OBBK9Lm4bo
IqOYp7eg8eyPo4pjzkbMGQYJjBj2InmltgbE6TzEWDjM2m3dWy7khGdB7RusWwaY
J3RttTXhq5xLMluj1LSUaq0t8U7D4hg3Cggl9WCKWIczSI3lJeGw4dToJd6lP0Zv
1ii647ZpwOlTPbqRLctqMn6YDrSSMJaC3twE3sUHTtmXrWOFsIguFVXl5SqAHPC+
+Z6zd1LNejAcYXzs4sNDHPaGoHoPS5ZmWUL8uvXEwCFUBdZDZkcPAPBTF4qhxi3n
wUKqE2gBetHIDkbcZRxK7fZmSBWAeEeJUiz70VDOugFI06sNP6KFDajjOF1Yuet2
Ikj7R1qMgrqp9/kb4bOEN60cifl9hukeITWIizNoM480Le9Ki4cFIUazALVZUr/f
1dwIMJDnhb8cWtJraIZIDrhKn4VvP0sLKNMN9TU4W59hj4Q6l+MBAPJMjHaKsvnu
gbWhwaFQVV+c1beDNG8wwLSv7eZZNY0bQ7Fe0n1VwZ7g50hDnQXsLv5eubUVfQcy
eb8rRKJZYX/mKTzBVVkeq5kGHowboBQewyM7zYGN7rOf2QRaPm4ooSwRZCElBmE2
ugLG3+1XcyTCDeHfBg0qh7FnIHlVyrFd/90jsMWvJOA2Wt9kStg7P/HDqSybtwVH
0y0CFyDoHxsgLisDbgzFri9OqHx+OtLlC5KmLQIgzYsTLL571TwKMdOaCLYUnzkq
pl5scMruwH7De30A0zRYtEkhrOTJ4um+tn2lAbO1JmA2BoDJT+roQaQ2Ts3xuX6y
`protect END_PROTECTED
