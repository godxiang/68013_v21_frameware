`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inmxkRIzwyM1tT929HkSpAoILGFEUdhloICe7e7iGZ5w7PPwc9gfNnq2l8f3HZXc
ioSDleGli/F960GFpViBQp4rhc4z+ZRF/UNDl8eARqCwivSygj9etOYhFOqqM5Dp
VN/2Rh4xQCmuwl6tDRCMdYJT/n+d4vR8MHGByYJZ3UA=
`protect END_PROTECTED
