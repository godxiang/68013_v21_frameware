`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlfZaQdsgJXKvn0L4abR6Pc0l+47CDGZ1Et9bUeCu13b9lm3wb9+LZHVbdcEMOrY
gqe/ep40NvOE1XjyuzOynFKyfdx//4/d1ywC0aLtl+6IKJtq1dpjqK5QvP5b+Qu7
RoOcHwn2eb+uGKdWACvht4Rc7+kdhIKRnxq/upTaK+ga1uMW5JKH6C90vYgWfx6D
CHaeCv3Cx/P6v51TY1zjIjGX9xaOgMPkK3hcly7lgMrZcmQWLJG4O0sqRtw3X0E3
ZArKIalhHi0ek9TZIT5gv/L8FRqW+jDWg9kRSW9SuSPhs9Zwx3VZqSFUdqxBgigG
wcG2Lokt6+NgGBTY1khVJqmhZ8D/sWj8xVuwUj53+Tz3ym3oKHrtJ5ezNa/C451d
4C1GhSPj6cCnYgKVbiqETHDcn2lOy3pSYnqrWtpEoR4Pj0HfWSDo9jdr7AekPUnK
tgyurxKm61SZBhmtmTZ/cXmaz5+equoxI0SzVEkX2Y8lA+34qn+KtgKXT4Ap8wUs
IXnPEo4k8Ma40XHpB6hk+r1fEcR0cq507rw2k569/6A9heG942B8PMzmOoJxIDnJ
MB/jLKL7+wdDcpwnWwhrMJmgNi21e/rmwuh5DkueK1JoTQ4VBvzb2HRrnCb7Knaw
bl2q3gjQV9QpJT7klS7UypzLTdyu87ppXPQnj/Yl15yaA/RCBiquEwtJxlOa3usR
FI7EFAhctfHX6nIic1uFOStS6+NgySHiF6HKJ8e4U95M+hKXX7XMoDnsHqEqslit
xnxACCW7feMIdm8TnptL9nYo2jBLWe+dSYUb9VRVAc7MeWL//tF3C1EFoafPsvTy
1OM8WJFV+1kriaIeMwFU3/4qDCEahj3+ZqYkxuIDQZIy8Z+0PCGX7/gnWu/L4AcU
u1CtR+pa28+PIPkHKLg5GOqeAOdN93kOXJfEtLLauxISZdsp0TND5wg3Tu9BIJIV
pxUBHpIbswAiFZW4iyLYQR0fyhi7fI/2xMeD1OuuV+RuaVGwtoWEISV4ogRGkp0S
UTIpVtF6bkBKPiNEi0O7gaMPsr3hxlZo2Ltm6OgiSfI8ETCEdZH9KvFRc/XRhEZo
pcXwWl9rm+raVUBiU1BO8zwCaZQ4VkPY1RnBFYrM3vcuBp9dyWI0wOaTVpE2RCXn
l/lf1MEj4fAJGtXVnWUZ9sIJhWOyD85Pl+tFus9s3rLe+eUSK8UC3i1gFKEDwW7I
vRqlNCylz+dgvecvK4ZY63J0OsMcBfwQnLLPRn4wet746dOgLRx6Clx3HU7nHqr1
XARHe5uEBhw2mn5xPipSwZI8sWGPpLVouzY0yPiSW3CxNd5M6TLxXGyE6QoRCjIp
oYaoI/yX7Y00CCj7EF6UD9tEd0vdWsgv6eGqgh7z853xtX0TSK8ndqi9cgKsDU4/
mp9E6kN4dolUxyBk5N0lgepAjQ1FPC8d0OV45q4I/nVkhRu/OjTIBOjtUauhP9ow
waYyMdBnarEspXl5RALsnddwGPIumJPD2c9BxHYmXPXQLiYR8rw+2lc/zQmfD0mB
2sUkY3e35+81Jz4VyaxpuVavEHcRm8inVRhQib2GkGiQThOA0v8MOOIOwxmBZa0Q
IlFDbHNcjQSEnK8LF7Am2WvQlncmzR5zlnRneGEeVvLJaFYH9KaLQf5uRCLb5q0o
NmsjRLjhMGXJnNsxp+MNLYGJYB+a6qMie2tQpP6EuBpH15yaA3ayZQ7xzCV60VC8
zu0TZDZWVPdgU3qTXsRxchUKns5oAzSRB9viRRDKsI6NoX9Ky2cHz5soOX1o9H+R
l0VDTc8oiWd82FEacwtrxJKbT6I4934LUTcUDN431v/JEn4Ts/1wh+STVKxkLXZQ
OmlXCGGbtHNiRlA0ovRa8H7YVy38Ubzf4YGlB7N9Bk/8PFtAKDM4+3oJQ8vp+XY9
TynuGezWZ/QOVIEuKRVPyAVqHCwtKGqMRKnYbwqAZoPjvp35jjwqOJlpA23LmASB
iKQ+feVTCdF8gE49zGuqsQ1sCs3G6/VXc1ktbkSFSJBEN6qZdwKYDRW5IThBf/ck
mCkrr593w6bg9PX/IOpEclIXPJ66knZ68vbMNP84WeqetHHM4vzHrBOVi50Gv8v3
NY1m5X2YhWnXZf0mq6Z4v9Dpaa/+nUtauZIHnIbxvX2Mmmbmk13zOn9DdZbsf8O2
YzP9LuWnIEc1Mf+FM7VEECH0dl1SfJ01nK9BU+kS3LSTCWRBD/2CoLCP31WQcjgw
XzVlJ4pZd3pR5SYxQMmryijf4kuw+cundq/hZlqzUQY6eaeG2OcYbZ4lSv6mRHyX
Db12+82c2tmOEaJQu9MKf8w9A5Jtak+zK6/l+gNBfzbsl7ZzHiAeuMjyPfHOx+O9
Vw60BtCkw1AVjcmbWcipV89d9hZxowHWVw3IlibUDw9M8nBdwJpLhmIvQvbEXtOK
jknIlYkyq9p4RrwCleR1F/xDnQt4L4c+tHc1cJWkFMuDOYiRhzQJjbz2zWG/liL3
HJiPqbd0PxyJlXWhC6Hse+f7eV7YyGwvCuxh2KSIRj25Md9P31eElED6dd1iqKkb
aVdVXBGZLkgp4vAWfPPBt0tLHYYrjFyV+o6QBCOQyJmRaJyH4ktr3mxdZ8CWM1n9
qSy6Wu7TIBFQ0Asvxfu+AdAVR+UHX5AQNqnaPtWqEhmtSi6vrabcYFGSqZP+81oE
fCVi8DM1RnR0AT2JcQGSA4ql7pEAfJ2kfHZCtIp3p9mxBZqU0ebBZyIa0sfi/zcX
1hiZy11qJL+zWcD31aFw0whOxhCbsPw6tF8W9plwPvbLMqgAiuxm0v1Ka5/zH5os
K8uYd4BjpTpEED/FJeudwtFaTBz9/FRpur9Jjd5uKZfFEdHwuYZMTD9Cz8LcqvQo
tuiDGBIdOdmxUfRQNxw7EJwZoM8kwAQz47qhEAeOLfnTyn+akbefYqQJfpCMUlMA
zaY94NxcRPVLXrAVgrb/C9y1yicLu/jV0DppmL8mm8JHq1+yBLsnHH/f4tEXBvLe
sLMaG98bDhFg80ADy4dXJwfgyJsgbsyt0aF90Iqa6+UCNE1H+uaMK28FM/bvJHXt
jthnEHdqTGw5T/Ilix18AfMbvAyRN9k5mN3T0LP0HslybDeFX1MAjQNfwWhWFGBt
I3+/IVbVkrFU+mwM16+dCXGSDlun0uSSFWk1LrohlMecLPr5EiDOn1OoiK0HbjtT
3d+jr5afeeDefjGhl9aUfuh9Lg7zi/0vvmXBQvWMWZJcdAwK3KmuzYV09y1zKbjE
BqHHIGH6ih8pqKsjl9p/Z8dcOby9JQx/wad8tMrUVbJUSLsWZ7236Y7esrIXpQsg
OJEtXGpiETbtfJFygifUF/z8jAii9O7hPgpnDzeDx5U+I22EOkL2U70+DSpB4J9M
RD85gB2Iwhde4yJnacgHEGa2rXcwLhgmuvtlezY7/92hkXpSQ6GqBdqmRrz/h47F
2JUz0GdqOGY9TU74AF3MTdV8KGgQaL0vaJLVuNeI7RT84GNYHDXZ5xCZj75em5I8
676p74Uly9o5e0MWMGZQ432PWwEWEJk1ZsDLPZ2T1AJcxX8TsBcFOHA4pD2uYBqO
iBtsmD6887ozFATuzUJud4JsWfqSAQLOLxtZE73fZqAUX0BY4pncST/uqqAXGJYI
Fc+g6jxbxX9jcAtmtasPyaJmIm0vnQMO+ZgnqjC5fyJaE/xa66psjnrFOd0H9Tt+
z6STeOO6y+FS7xszdWIBFE//1n63U9um/PqmYAKG+7GWYQ731v/9CO1OSfz5tiJE
zA0B+PjYbSFy5l6Xap55QBZoidKULhlq70KdUFXcfbdCSSYnSISVEOVK0E+Wtwhz
X4EEtNsu70lj6SCzW6nBN3TGafAOfQyphsHn936QF4+30BecVQbvFsjpW4uGC5zH
zpr3HFoCnikaFmCmTsO2TyW9yGAUAd+bsJGhmK1F09hOwbXQA0YpYtNF2tHcjMh5
wXGpvsK4Ps3lk1N0epBsXMmn6YqDgMNFzIOJbqR9CLENp7/PIFowkbc7uzeMqWIo
oFTkAGAuI+RxW9aOKpWPqSAmUOKw4JOSPCz7RGln+3PCEeEbTExGtGffKCICngyP
U350NeH9M26XbsceS1NtiPUZ6YRylNa3Zi4op7hpdmAPMHG+cLwo8sahgZfS9/R2
0rbTgCTJ77G14x7iaXtfEGHl+G0/ntSAQ1l5hvN7coMpihKdqOknpL8T31tsnKmd
tT7Ie/8fjUPWJFdkm1U1QdKEV1TrsgGLeQHiqKHI6yuX/Zo/hGZFz0PciyGh8kFo
k/shbH0l8XHfLNuBMj0kyHyzoB+GDUB6zL/myRHKQw7EP2gvcEEi1oqy0kzXvkde
N4v2gt9GESLIAX7jXnBrDushVhexrHdJntcQmBtkgcSvvojlMgUcP/OelayRDtZb
pemQhuY8Qds+9Ssdd2ht7CcCWhxM2UZ5lFBRgD3ANuE059H/UD8CjbXHhLEoEyph
xToB+v312i4lroaYZkvNoihj4tEIL8jFAGqqLNE8jIGIHJgVOCSmE67hEt9GHBhs
uPXHDfy2Lrgo50BbBGqU6rtSetr/cJIy+4S+XNt/N8sozXcNPOLJauZUYTdtZ34F
AlrVZS2xV/Eh6BEL/C0TvUlUZEcl9NT+8kVaBFNqfjhr/vLmXId4v0DpuQ2ykcjJ
wuLcfuPiLpPvqOKJHCB4+e8X4PHeQf+TKywawKkC1tggsBZ67NfTIeCJm2F/qi8e
gcNlS5iw1XQING+2e3V0N9rN7oK7640CmrEwQU8TtJTy95k6d6c1LBfd4WjXX7UC
KI2pEQjT7YSdTbW3mCG7FvQOa39xlWA396rI62vLVGbZEQX4o9rILwbWwVmm3wQ9
+gJyxdzNkxGnZcEJrhD74CQzn1UC3Bwtjz+8G420cbXK9Vdvvjzf9kwmvMjWS880
Hc93Z6PqOIb6X7QgIWXz8Jh6lRW3PGvVuMW1B8SQ9tc3e2LeWLWCfs6DPmZ0jZFU
ChDcHEIRg1z8qHC030XhdB6JhHQrnBsfW3FnJjCez278KJ5sDgtTF+dxt4pnvWiv
2DFWjHhSQ+cdOkO76aR2aTKKv9pQvOMlHX8NZ81Zv/qzNWd20eYasaLNpdnWg3EQ
8OCF7hzJX6trfMgJ7/3lDlzrfS8UQsIDLKlWvdRx1qGqfolskexDNvXzvvdqXYtx
FpkMdVu896QGMzC+fc9ExNEz5UaCfZzVfwR3zst+dwat/lqQgxESk4uK/hIrfEog
+IjFDbo3XC7J74flOh2/JPDYtq+CdEBAOJC3VU5ETgOXLAGlooyAI+sJQZzqq1P7
cUMmFD/NaAtadm/YOO4NliezBakY/HX1aeviHQ1pdOap+pIIiRLXoAnA+o/JDq6q
T0udO1gH7AwcxPL6nmEbed0siQP2lxT09+7c5UuWfXW28Tn42ksKsta8purwbZDB
UxEo/L/tEgGAHeL80jkDqVJeQDiB/CgkYLkfB5aob9LKTONji3lxYkmEy+L/GiB8
6SDzItw6rPbZn3N99jj28/ejDcoVvcu2SeSaQ1H+96e/iZv+42Fsazfs8gyCeNRu
qNfQoX1pNm4W8MAj+A0oAwTghDxj5Uq4ciwSvCcVwMXzZfw/3YiwfEoF3bJVgBpu
CnmI9GsipXha2gEB25Jn08NIJZS3Xm9qvLobN8qWihePX+WIs9YWMHev3pmQYcMl
XLKvsh6szPSWt2gdPM3Lyq9jh+5W2kbYS4kQY8cerjSpuguLye16Km8mWeHG27iX
M0+HXv7HA/IpvStDnvfM+BvcEylc9HE2NcJ+LT4rstQHHi2LItakS/Lb0Rq23Hdg
YNcOO9NFWVnKbcyBQedgVfd1sPbxwCMP/DxsLHYzjM5TPuJc1IIhMz0ugzVhei5g
fRGhkWAkRZ/+Yn/ECIYtBIvX7ujbqIpbdI1+Q+Ku7r7BYwfkJ6i5hQkmKVPXrAXa
8TOI/V8VYw2ui6gIDAih7cEjNxRnGP1sb6hDCV/262srn8c3XZyaGEe5imjms03d
eof+2eDys/PctEwJKaUKmuKu84/4p4Hj/IXd6c+o7Coh7Zt22vEyzLZGmj/LkUEM
Mo8ihnwSOAg1ZldlhDWqUadPyQxd52UDyVy0R3sBR4boav/gMaoVb4AyLXp6lWLF
Jz4plFezIFnL57+K4mJMZaVjWBbbZUoykAx43Pv87PofPB+gKKNFRAZXJ2ByGeyM
ejX6eXgK3oBvxS6yzWzeRpIDpfIST295TI8yCJimP66O+M67P/D6p1UEufD1zGwd
ugU8HN7e7jUjPo+tc6aTyNdxHjHqnBwcJq0rLydofh1HCpYBUmQT2am7ZcYD8/76
mAlpx2K3tIx43GQbJ8KgtzH+kj852mrFc15klPA16wopsCTslYVe4V+6/sG0YGGF
kw90C0n3ME6MOgS1BiUfLzF2IOaGDUkhfmu03jwkX33Cj3Sb0bg2snt2ioz/pODF
bF26yM9bq4vaHTlUoDG3MAML2KcbigtXSWQyT8gisAg4fdrBMC7eQlkaC8RRGW70
hWvK+KiKDZ/3SqNqsXgnqr86ckqlnNlcqw2YwAfYGdqgmtfqW2DbSXCJn8D20CuA
9OM9SC3SzQvSlmi3vU499NBH1iRKtHo0zJ4nKogyurgi+0JWB+/3VYDh3HLUsheX
L+hH+AT0LzzEZ1XhLu9NODnpBdVW76B9ebs4jNBtkS5nKIFeXavJUx87BXY89hJj
N0xrEWI6LRKCsuiTLHqmbm27bK6T79oqobNC02xItJ0+hP62d6rkNEA6A10E4N/x
Zuzjz8c+L8xp1YhFY8RDv5EB7cWBno5o7ExH66oid1rgHmSpVLNQY5aCFIaRssV2
Y5bD6QLDEzKwptBZqlePFqIe+DxYpQWLkQFfIqnoRb7A/xdMm8vZiD1rk1oZDgDX
UHGykGisfFX+SMZLHshXPrCzox2FXz3EFsvwgc0SEeCMEZGJCBO1K6LX4pePnzWA
kHj7dd2Bs1l9cVcJ/0BKAHbLD/0sCjk1twlYwCM4P6fv9sOWvtm8TH0gi4rfOrmm
0yaR1CnJ+fPmm2gfPe2VozX4I5Mf2bAMhYNhbLDr5aneOT2fe6CeiBqS4CeP+db+
XnUdR5Hus9mtd4i5kHs0tcJD9kFdDjZIx7uWW/0/GjWZlnOF35y6pl0N9O9ghi1a
MjKG+kFUMzpU/AGf82ac0fEB/+JK+l3R6hAW1KV3pFCqHVvRMc8CyR3a4TXhmhS6
vSDyL8LaldXAECseDQps/VSuiY70X3XbSopedVSfuSy/W//k/qKbvhxQ2vn8PfOf
z0zqDXfBHOs65dnnt6qFmw==
`protect END_PROTECTED
