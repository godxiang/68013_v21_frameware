`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwCsQbGerdqr+fjopzbdQq2CjHXYAqI6YO4urOqNnK70nPbQDb16w8uvAyUlo7lu
xV8Yazg+1RQKdtMozgK08MbcSxUKXItThEaeUEJBLZpa3Z/jluNpc1MkHHVvcjEa
Dr1MUXsWrcW5q9OlVzAmqeqrLFJxLL68xtm9wNegW+ryajkYBcjDZfd/fjYF2iBg
WAQMW9cvqBQDGGB0OmAdKIVIGWhlsTe5YrcMcrZ6YgeZGLk++IOpRg9/vRuV4s3M
4WQP1evx7x+iVSbCJZuDp3/FHVPZGRolIVb6II1KqWU4J2xu51Hjz4pz2GCulniS
vEypBgLJSaTd03YzLQ2rgn3CF+Uo2cwzsSkA/oTqwS+eVVtByUT9ReSqM753t3GZ
KsSicP5A/9uCDxN13fUb1nBaFCSw3EWeQES2ttMv9ZihKIX7EbZ36JPh1OYKPYdV
5n4N4AcFR6WryKEwswC9dmgSOtz7cYpzB42yEpgcyE5b1UcKIteE3CeYDymz0O+q
i+n4pmhZCl1HGqQy5gaiAB/8dHaEafxcs3JkqOppfVi4ko1o/Bf4FpyKW7OppsZO
hKlo5bSwGhwuZbRLHmYpSCY/DYYafCLOhV/OrVwi86VliWEl4wWSMSHvyDPca1RT
ozpErAu06CxfpjVuhSuSdy63yY9HggVMVttewVjlJTPp4PMlKPVRYbaWALtGJGHf
NNGVGW/jZji1Wg8oYbN6yePLtXQo1d2AHwJHwS2WMnW0FKDfHRxbo5tQoLQOldTs
knlPFKI62LfZ0cx6dFHhhrhLwRyYsYt/n6jtGSIvaN0tHX4xX0fs6sjDgumyI45/
rteLSQoRGfTnYT7IAjDaXJ1XZIzyJnc+txRC/+fsLDQaa5z5Yo83takLsQlMjAV7
C2OU3tZKK27RhzAYj6ydT8IigloBFpoGbfSzJ+aETtbR3rAn3UjRPbIzT6Nv6w9V
XNZojsyeXRSgPG4NXN1no2CZTUOAJVbYABQ6WX/7RciOFmzSsAWMk9uVBay1pftw
RS3aJEadMq4JxDvdAVKuc2LPzfpvL/8f2fy8BeGVVHdere2qRNar0un6/gsEJA3L
84qZNZJJFl6w5KquIDfbOaeUwkjy/b/d2gIfEf9R5KQYolW/RPN2hYerLYYWjBDl
xohmGslbt1WH9YjMo/cKFriP+XKK1zTN85SRtp1aw6asG9z38aQ4KV5APFN0ZPEo
4GNgjsNncYUGPgWyp1SFRrmhGfgMSsfMNeDR2cm79CU2RnsqqK7u/w5MbXB/1Oor
Vzt1nLsBM8BTRDvpKN+kcPjX7kTugawusKeJ7wUvL5J7aKrP4ArHMoDvSF5N2xac
eNEhDRBblSdkC++My08cubkLbXnXlDXA4xkZNvydkM2luxf9GT9tnOX5uWtqUXKB
vekwPvozlehZD4Qk2Oujka1Jlq6//WZGuyYSS5+0wD+fYA1RXa1RjWNYUiI8AjjI
dmRHBy7bSKpMHOMe8aWoRS5p3gHHckMnjJAzyoLZMvh5OdHZTUSd1RyXjW1vVyLb
8l9n08ESKVR/laZ4DW5aXJv/D8un3iJ/vEpKkB2X06TkQ3bjx/lAEhLTEmXhwEIt
IYWomiUOdc04Xv+/At2YZ2rv4czQ3bSJjFCoLsjrljwQSluUwusTFBEYnXBAjD1g
uHGOPFcoTG4ssQVDh65L6VuNPIKMYFTv36OiJoMm3sn4NLHQDOMbLSOYq2JFP4Mn
MowlRvluuFeByFRFKK4Rw12Sk8LiVjS5/u3FtZ9izXHqxdleCdNTpSMVxmAvVZMj
QKoUtBNn/W9aWuDp9EuzRLcDq5szFKjt86a5+CaJ43yeDnyavxe5Wpskbf0mWNgO
+UJSAO1KDR9IUcfAVtOjyinHxfL1+AF3x9ma/jCwy+wrqOfgTCO+SP+taxtAiKhz
WfjNWiFHqZE/nND8Fcv57yikdBSCoEG5zEEBbs477+2oMA2gcgj8gJODcTtmGNKP
zTtyjPkgJDyrZljqUfIoY/xLKHpFDRybHWAYO6PwGK7cEJ/9f4D6wxAThzxlFEH9
WzW99/TrujIY76GPM9pWJsjWQSyb9v2dJ31t2Pxf24ISMaPGTEHhLgpeypdkrFbY
eVJj4adI4RicpYsAMeo3D9+JN/3qiNgKl9EwgRnayaFTz0JkBqs7aZdvZFyUuy16
XowSqLb6clTCvScsWhR6Xd+xt4nkw3blyTIs/KY8GP153kyx0/Q8Z+DAU4AnTabC
o+N43iwwENgi01viHeq2AyQ/Ts5zQyF/SXy12eWIIPoxZr7pDaGSkZGwMcV5i0bq
OofgLhEENQ5vb5vEb++cnwrXObhUlsPbif8yo2N/wwxRIV9P5KYu949rE/HQC80m
kyiK8fiHwuBigkq/pyd84QmiWFDUn66QrG7DoQr421KLaWZAoJO3Gi2xZP878C9V
sOLODShrmBES6pH6lGosjGdbxa7uw8LGvd+0de9ih6uXTFC5u3B16zZ5yBj3mzNr
RZ6pP2QM1a+CBycACZdC33pvCik0iLCTPW6TM2LPUXj1gFdwkFc9RYKphfJ6WWDE
xOE53kwT2ND6uayyxpJp/raMhLogoAFAbEuHDs8hmXF9PALncWqczwhYjKT4vSRf
h7C1RtgDrtrKh+ZlPZoDe9cDHzWJkjGt0RhOMtlBmA5ftMgyfZ5UCZpXiklK9q+A
TVw3gzim9tg5kxmmgBHAFHAlRaNNEJazk7cDRpjXce1dNV6fcliXxu3LWpM6JB+j
S8/JFRpnkKeyuu/MNU/VwgGjV33fydcFu626OlFytjCS+wEAT3zZVWmcXeO/7zTo
IkMLPYt+o9z80r4GAZQ7zohbC9lGzEckVjRSz/ci8LwCABZy0CRFEzkEkED6SW8f
yAE0OHDfXaU6bB7LPK9hsq2xB31H5Y7DHl9Q/g9Q3s/edXei9RxGQBcv90/SNqul
L5rYJdvLratKi5z4dzec3yAAmG1YkctydrVmUUc4cgJHq9igbZY2rY/5t7HkwcQ2
NxUGaSS7Buyk2gOPB8jt7zJA9qDy8pS7g8LriyfRFqLlm/zEMwxW77shtVHQ3T6z
ZmGAZzPagMwcekHh/uzMdR1uZ7vp5ADRz2d+hGn+XMesKbzE/wdmYn8l4IvQ0RtG
gMJMoa9IU3SSby22XnaZgnyQzMGoEUf3Zt5z5qx2+oBdSSAT6+tFVzs/hXhtyXLf
f2el9NAgvjHyPmt+4Hl3VbHoJsCTzMrf+oxpAUwvGwntbkSl1GkLHuUf0XoCHpFG
etbAl1g8TWmqYIY+UzmJFf2O2xW6QM/c7i/QD2GVQUhcbY5+aG8Aenj0nhP1L0BA
EU3ytL5gzRQyUHfHzGyeUofaBExFf3dBlCiUkJ/2pY3lDmvsOYrclJvWMB5yc9IG
SFpa9Mirp5baDOgfu60pkuZSKMSu7VGX9gRffDU3NosfVRDtFRgcoLbSRun7lWYF
2/LPdKS7QOurbArNNEvjBn1EwNAODOdFFjDs9RmgpjWF6BspQS8kfZibyfvfyI4l
ZYv0+h+LSjnvfsMoD4kfOSfpvZsndMAqvy4VYYYa6Ct8+ek9SKnd3Thuhyf6u0Hb
We4K1+89MLR0tYzwYfYAwuqEWCDikVlmoSLbQ+yNlZ/0mIGjOaxHaFmKm4/WS3NA
BYYP2RCdfqD08km45fEfCpGjomSbZNFmkOqje46806fgIj58eRwkfXuTXeFsMsJw
OUi/vENDd0IzepL4E6Q7XU5l3o2P+cUkCZ8CTBKlJzuNAcj3M8ZqHQ1JVUJa8+BX
LZetvhXGZLsOBexoqE6ZC1JHi+FqKxpV2kn2yyJQCFbYdoPURzR8nk+u4lq9o5WL
FR/W99BzsegTDXBKWjg/dEeVVov4q1bcYr7K9IxUXHcRJ9fodiBsRHqVnUdXwvYI
X00hF1dYOjH7oceZ1vZ3Wis5foFg6di86rqa7jkt50IoXh25jMresF1UWtB8UwA6
k2Vt8XSyCqEo5DXJZHHUYlPMmiJg43B9eNY+8BJtbMTAsMFKjRCY4x5M7MAe76Zs
R+Y4VbISuGpTULMrNKeEQ4ONEo/Nv8Rz61xL8x0C8JfLMggFZlxZLfj0iEYUVKZF
5m9Cc/gkRzkSc3lM0d5eoUt79s+uG6hixaisYwY5h+QbhZBKt/TCp/Pf1gEeCtfQ
t8ILYyycvv+gYv7pcJwSzUV3XGhn6Ipx5dLOgKLTgjQAN03haNehiNoNrRPZtUI2
LbLsoXXNpezoaZK6uH0tXf2iFdlqnRwIhtSmRI92fBMcTiGI4mmIxMhCJJNvvfIs
JoNJU1R1seRsyoYszSws059qWXoXKYN4AelFl8jqJjdBfRtimlXm6GYllnzL1yMq
IuEWbxd+obAq3GcM7tYMI0TWLdF5xhMRNeFBBaZhfTXTI72VcNmRYHXp/NFKHObH
MtWJ1Sx70EL+oq/JjUuM8RBlvPVhoDXjuuLWo/kR1f4RLiiAy8VlYh/fbc0N13Cc
4Rv/8E+ENVQVxuMNdPx3JT7mzSC4NaNdhNGNTqhShDayA0tyT4x8insG++lZ/nr7
YHbMoWaAZGX1x352HlZAplQ5FEi3Qv2KHqIMh+qQAYQbX7F3Fd2IwY040ir0djBT
yYdUsdh+ZAcgLu0tAAOQssx79nAMSnYrdIe8CSJoj/2s1PtWyFCdfSyNL4O1yI+c
+G391VjQKPzlXpkIusT/KI3X67NeGgwbEN2fGQOjQI81zijOaims5ldHU4T2fgIa
l4Cq7fbTxJInvQHn4QeIkYRLfLxaGdsFk2Ah2ypqBaYBbV0uPtfHw5Yzwx6jj3q9
zzwaKSJN3Bm+Ha/Zo8b3/GVMaEu4dE7fLFVV/PpuF4XFW8cJZ/jvrdXFbqc7vNcr
wYVdglaef67tzqlC5s+n3x05BwObHfcwYKEn5ZWPOnAk8o8T1beYiYZ2gDlbfrPN
KJgltZg6EiV/MOYcMXvXw6nS0aYyIvPmki2uV4tICo8gqs1YUmOJilmUDo2D0nQL
7Q5GUhjCNQeWnj5vCB7J/FuE1SSaNNDfyUg4KWWNnbXuIE0ONTu+d0CG3UAs4kXZ
0O3tjIEV8DAEOkinR6yFNKjhAKwVNkGMkKLQZoCmyS0XQ+RTw8yjALFXcPrAQxbh
IyoryItESG962IEoiQ1D+ifzSDkRjUQeIJsGiku+6B3AFdI+ML4Y8LplnFl7S9JJ
NP+MJnd/AN2WsyUXl/XeKSimxQeTqFAEZqqyRQev0RcFuW5nvlL+VGd67iAuRBDb
4ubquqzMLVDtVQztdeKy1lLkPlrLc02WKdhSNAZLx3TNEIq7gmdUz/BQvtjeU3K2
GoeXd2aSP0TiQNJ/z/QdsvEyMooe5xH8tQJ5WdLV94tDtVMah7Wy81XJQ/PizthP
QwfeERR1vGoW79hOQbESYle88+3k2/cKfoeXQwxUOkKes4+4fVldGx/KnHEuuxZa
X1KQgUSTgNwWMsTR9PJrt2q0R9RkMMFVDkRigtosNeKKDL/uLKEjvAwgm7AFb8fY
n1XlX2WoLyfaCxJ+eyTbnvOukjosr3iRAxoq7VFNoybRFJToY8GBK7BNvVahHaj5
gZmRjEnxONoIljKC/sEGGEpqkhmceFrnvPlIX3QvlLDhY59SQi9+yCZ5oDUV38Mr
bZqUgE5Cc9H6rm8y5aQCYGMjDqcKx+Odca7yrJmsgmWraUaUVN+ieO2bf2AdRBKn
Y9wZxdZJygo/L0vWHy9/Kg7buVk7kNc1Rre4dN2c4LfeH7CKOuh/r/oBFa4Wjf3z
lEDEPgag+DpkMwVxgPt6rIMSnotms1ELrmAnBZ1VVuMdD0hwm9XloFhl/Wo/kicz
wYNy47pG1mSIXdtyZMK7ifL0at0qqQhuBTl++HiwFQRp6Im9REED4hd3KZwAIE+l
iEUC7wzYtiDldVQQ/AslhQ0i7If8ffbYOWppCvAhZI2MqKrxZmdp6nNPOnwmKo97
WMmaekb4BE5zwtpHNmoXlsYhXBaYn3hNILPzmrTWtabjI4m/WQsTrn+IBa13+MN5
qBLfdSRCXkzxC8Xwu1CVO4wbIkARHMrZKQlq+VErFuM2FesjCvU7qWY6aZ86ydhQ
WKeeiNdqBTIQYgk/M+V4/5XFW4pZypeFSAA+LoO4d7YGvVNlcsxiuMQzloLxPqp+
I+qVUjMtYxr6fxxNSA3mO7ToJc/aE+cp7PanwQd9pthttDb1YOuZRiro8sQKAPgJ
5znwKY/P3cpXoIFspjlZohv28aHaUxImG40VO3UwtC7/UuSFTCLIV0Hdq6TVkbUI
44l32fCp3bkPKb1vZFuhEZ3q1OEucrNc0f//w51tWEJKdENNVNomRNwRc3mqTmEw
1QNbUISPFgBzYQGHLTshnq7YzeNojud/kSA+OITk5zPTxGKz1ch6bxBuE0vk1f2k
25KOm+NaAyS9uTVssUIGYoyAp3478NpDncrRW/O3WFxSO1a4oHaqQhDpuVxVF3Kc
rH3iCSQmJC0KlnePljBIuqGJfou8sIys0D7VgQMHIBtr4f2q7Hx0RiK7GkcHeBRz
b0/QgDsXt6cJWCVSGzz0RTkRCT5535B50hTxvw50HLG9BHn4covMakQxvZ8a6sjP
ZcS9YmLVwxLzP5UwgnvgXmZbHERgecl2wMqyzSAVRgJ1zbEvDdWx4uwBDVs4TKDx
baXwZTMG7Nkz3MK/edOkZaU6v/G13ROJHzTGRfIU+SvFrt9AF1Ynp4AqxiC9fmMb
kl4Wb5e/r9jNcmt6LXaa3fHTqmeLhm4QE+FdfJSgmGswPgtLXzqEKbg4F7+Y6Fyq
vFsABFYAGU5N8jp9h/FhTK5H41HfsMvPEQyzpmotokPlA62PxsH9nWYiyIYLs3T/
32HQcHgdnFqfVXtfv/jYlTLkduRxAvDr3MoDgFOaYkwyjLlS4ZWPhqvqlV2O8HxS
UGJPna4nx+yu8iOrEVuJZJyzGz7GnFWYiuzGgYfeEpSD37+t+Kio4uHAmIGPEJCt
IvjfNX6rY4uNCUyWaGPpJIba103ScZAUDKiT7PevWbRGVo27tjuNXsAUu/UPJKn+
iiIKT0gU+ze/h+9nYEsH45BlleZ1gRKDgMAfRf3Nl8LO5pzkNO3q9ZlqND6iUD19
CqfLa4FsHRGdgbyRBgRul/lvVl1XO+FttNBB0C07uZSXElYMyJKIeGemC8ehBGCU
DgabWUuetKzyJqX/CW46lqC1MQRKYDkKDXUJCcZZZp8oExgGzloEAeiDd94uKF+Q
bPdeG+PVX17eh9kSRhrJ8kauMVFAGV0pNpppICxJtM8icLRonaKdiHRybD/WmR6U
HrQGs2+tqQcjnRBqr2GMtAx90a2RpBdVGQX9uslhBVdZg35QUjrPk/1LBuUyceuK
ecDfTYnWJN2lecYdn+IdPo0WdGwyPAKL1pN9rxbNuFg3zd4ooI7QkwtF01+mU+B2
91uk6SyNAnEIy96GJUT+xXWst3oWAP3YMYW0dEdwPXcWr40fEb9CaKEGUzA3zOL3
cXoCIwfnxn5dj1knDWeKU+orXaMMPXuabzvqlJS6ZV9dNyNRRKGR+n9qfFlQY8qW
0n12j3XdNxKb0FV1wXHogPuHih7gBHJobeC4K/UCbzBr+7edOhGDsu686gCaYkLB
/IXbc3PbY2UPk6a2Y9La7M3fPqUl3ZZwtGfrTp0UnZwU2bqQgCX0sTJIe66jLTac
oQdJEfzQYKsuYMFBCDAedf0ViictAiHw0Y5FQL1l78OZiohQZdjl5NbNbPZ3tEvx
umka4O/p1ooyyjOSVDC9avD+XcrTqIqWdGQgt3gdggwHQR4zJ6d3EQPj+k02qpkX
C7EQTudA011XuceNsDR4AyHS3vCqaQquivlgG33kd36lPdY+zdGtmKVbOl8q3uVl
tG23/wjZ971kFSmwel1XLSqWSXojpwFT8qA1ue5iOQJYrD5sa1sQaPszU7j7Ca8k
UY//dIE5xRLR1LFakm2KoNMGqNwXtV8vIDeLo823J4U++OWV6ZKpfJRfjXw/egFU
bHT/+sLbBUdCVcawezTrg26k0eDwprpYVyLG6CG90IJFRJas81finXvoOFNVQY1J
Q1zbcShtDyDvWNSXg25khrXQpj/ucoID5xL5DPzx3R2M8Is0j2i/afZdAhCi6S+G
3p2cMETzkXFtGJmF8ho3VQkjzAOoHaqagjtDwszLukAjUNTc5S0P5OXMXCoR+deu
U3vp0vIbVooMiwmMnVVNN3Gg/tahQ1TszqCGJCZQ2inBREUaR7FZnxhniyBCMy7B
r7ES0Z2Ii6ZvIrFTou1YHM/R8Qu99U0pixjnEGHetKb6x3VG9YgMdY406xvCH/4t
qs1A7QUyVY9kJd7NJWRgHI8UhEmitn5g+mLbkUd6tftU0SA2F2LFBp7MRxWPtCPY
TMUroTWtTcZuAVm4CX+DwUF6DNVzLGPIVDBuiAbefTO8gYGW5j3jBLrKC1WNfpTb
bL4PRnYFqac6mmQzCtXKamqArrIk+6oKi2/pNw++8LwlowVK30IVtmbIEH0UBG2j
QOA1+PLlGKaUFEVEI9RXZd2Atbr3G9C88k1lIhFBJodjebqPIeiXzhaYnIgdhIpR
MOEmvPuZMbYxVNPSlXxXJec9vlZCdYU/35Bj4cgd9PZ2yxWf6ToBePIEFZJukPfa
wOfQLA/r0PWn9rGk6Ry666/iAVY/SX2Nk3/1NypD0H3ly35aTjwdZABQ6DkCoF+w
xe1spE5cm5RlWLkAjSjSJ829B7zd8NZXtWb0xkdaefNdef7aYpfdPl/v3kQVrM0H
PJdclKGtdpTpUC3CWTC4PVpNTpPnhGZsG/2Fx1i/0kpj+eK8vbK4v6d3OWT9tSMw
pI0R8ZNvkuWphx3Xvj5kmEXkJqwIzcPgGgKwUIZXxwVNhhbnRzZHVdraRgc3cfwL
liTI+zfPkbXgMARZLuyVEc7n6AOGyh0UIg5TbcvCvBwLNUbGsictYnfgK3Hryumn
nKRJSPM9mef85R96Rz8vk74LEC2AeqKsMAC3jx833C6qObTrx1E4ptjgi+kYxXxO
0F9Lx4LFSphtjJY0nFHCJvH5Ja2mjuLzd2uFQgEdJej92a+uMRObsXrPPt+nn9WC
VoCJJrpTVJTft81YTe2Iy4049P/59mvRaQjUtsO4bJwMLlqcK/fmnK6Hm5JzQCEM
ClpIqQPrna7Ta44DVj/P5fsjgHcZhbfiZbB/Z29VWJ0w0SVeVlMRLeZdr2P431y3
QRegQcWRaTOf55Sy5FCQvpEm3VuxjQNM+nkPqTVRs1BZ3kXLTBlPWrEitNbqN5A9
F5w7R/hYlnEzZkFcE7iuF1IZTSGN0c2QIoePGfRmI0rzrOJ3cSKkzIzuW3292SXw
Bvhym32DtXDRlQSKcUBTuBnjMlf4Ap7ntEJtlkRBS4F40SmoYu4F5onEHsMtfR21
UczL+ySoq6M1ir8/Z8mpyLdVucUh3K4m6DpQ8vDRS0UG/lDE7mOiYaUyXHFQR6vV
F+BZAG0WphEUAKBWrifkp1gl88W4MM7exouxH9dZzGrhFaR31oA8CnRfmXd49c4I
KAj5R1nG6pu7G1mXD+3uS5YfAOG9vSt+kuNMJqcgRbdhTSyyxfHM4z6+Tp1GQkaF
5Y6N1GomWgzJiaYmFMFb8J9jxUcwM13LibKbLnPUrABgJ46/8qu8AXmgxkH8MqfO
/XMzXdeIjHlS+VIcm6+ls3Q8MP8Zzg56tsdHy8AowM2zjQf3uKWzYd+Kadr50AQk
+jEXaWFBH94JyHjzRif9XDYW07u2JwB92xc8vfgtqZpw19Sb/EDC24ZtvP/XENKf
LX4OdIvXubAX2jbEWgVoC7YbIJxjPBxlri2qISi8+Q10wf0UkpY/9GFG18Nic0Tq
GIs4z26r7D2VXaNXxLTlIkA+CPmqhz0MucpaSzsL9KKpYzpPCtenMqwL6QJj7T3e
p+lGoO8babkY5x6+4Uj2Jm5lJExmDhwRR4qxV4Kt5qiRXs+f+44uQfilihJfsXsd
noZivI3ORIHteOD7L1WaAM0j96+sAxQTOLFDU9mgzdB/Kw06CiBaRhkmeutGdNvo
CpVaRy4zghg7GM/8+7rHvedGdwnFFRUlVUEm5eEyZJKRis3KXgPqzpNsWSPKzNMC
JiWqLQY1N/oz5MEVq2qzqxxqrmFn4wfHKQPpb8lzPOVV1JNmN4Rpg+09hGhHN9UW
s4uclvMl2WTaH3Bn4m6Y0GcWKXqIU9SspYDCv/VQsKJbLpRnOSFWXFQp/53hnJV2
GdDUMXV6H2qWJcia4gqVf2lR2XavSd0LHyHrNsnlC3KSXUkFmfpjbcImcUAUOAMy
8EC9obxLUo+RCH5IGmuADYvBKTycr12TWEHWClJbNpCspsBSqyAQjjgpu05aHoSf
WO6iiZw7+s0bRv0poFbY7n+SDs3Ir6KZP3SCcsNEzqaZvlGis89ZJ9JXjUGgZEnZ
2yGoCH2tVYZN5UMhFOpXX6gBkeasHE5MM66MZDTes7pL6sMeXz8N2Z5yyPPg+Emj
jiR6xBeyCQ6nnJf6kRTJQv8WWyYdb1lL4sdIEZ5O2+kTjdGb/vjkeg3egGdxhQh3
HBgUivjJjxmW/TYusoQMfOmxWPi3e3FtFhCAeryG73bS2Qf67RxUU+QRVbYfwEJE
8IUasOUvNKcFL94xsBe2JMJOgmIBJfDpC9oIdpUFLjMxVB08yTEINelrGiXArZ4s
ksCgPUAdYYHLDGuz7w0uKZxT02vhCNdew8txuMvJn8OPaaRxfUBdfI8Y61kd6A7y
Zor4x/rIw4UbU55c+jovWCYcQsk1JvA7zp/y0fQtrW4QqrEJDfYQGqAeGESQiKY+
Vzb0gYKxEApqxb+NkB6aNkNiy4E6VeCl4TS/THTuX09W9ZgL9rkNDqQDy1jriwWT
Xh01HfLNdf8+5WJS9AQO8CILKEOb7CfacybQXkAu4ReFxMjCG3cKoO+5fPE1MACG
r94o1Ar6+F1Muilc7dBCREdB1lW7nEsVJ4sBF+ghskapB4eNFR6rLB/3citYlkhY
SV7jHrlkWPQ5a9bubogNO/JAN025zIq2UNyovSXT/cJEBA8gIt3MK/4nhwQPNzET
Th74hh4ByIHByAxP+s7unsKewv4xrvAmdKRV91A2ziaym7xniHnIyrGJLdAJeZUW
JhKBUyboflLYawMyCYXpZgg/fdrMdKgkxWJyoL2a1kMXq1r2yiCqIu4nZ0tCaIlW
c7SUUdy7OP3pifQn7jGIc7NY6KA0dQLGWTlhE7jCtAAd7YKq/evTf4LU+BiDtEXt
7lr7M7r9i17XK0wu6y3QVQ0Vwai3AD5KYF7bE04YyCj57p2D8vBxV/mGqx5uIViG
HoJUw+y2Ep5GMW00b6CrlF32N+PS+gD+sjnlbk185lSHvi8s+l74wA7JOg3A9AuY
ErZim92ik+L6jeADL2Pyc7V08mOnsOmycVci5liK6/rXLtVNlXmv85gGFTYOfoPc
iaHY9wx/YRp+vvs080cV3Q/ip2XcuK7bK6DZqK8VNSkLK2SoH9VgRHOA3L+DIEzb
bov1QMenWwP6HErKUW6KOjtEICglVSVcbUwadS18UUmCr2FPJSYZ55iAN3imzF4C
tS8kqpvD7IeMY+HRTiIpja9GeKGo06qN0Np9sK8LO96zHCXGnkR26wdk77h4Vbb1
O4doNfk7C+eQEdjXpCGbPmN1h+UDA7zBx+91bcK5L+hqTCF5VxgKev7JPVswRhPU
7IwHBmP3c/YPP6RPry+maMhZxJhZ1+/ufXA1mQo7BiQ/fcmy0T5PQszVC08D9EGh
mv/Tj3fT5SvXXT2I4LSvUYYOhAImIpFwUKLNLEkKYlwzJt7TT1uWMLMrMZWKIIpf
Lmrte1zMvwwDBEvGgURjvVZui7T6d6mouZWpJGQBewxmM//BE4Sg9QZAYKqv1tMY
aV4s0BM4McksTSQL52RxP4fM28tQjEc1EacnMtcnyRBITMtM+czSBPdQEZIANTwK
ovjJLCYgAxr+6VcS2dUKRwuT/J8Pcqa2x2P8vBj+XVRA6ItgY65PEGEII1sdY90c
lsnZ3wOBH4D6WKh/pihYXSB6aLwrnp4k4Q2UBiDFr2z7PWmEeGx9uvhQ/Q5aV59C
rGiRH2/8WFCZ87BTZxtKU4Kc3ZJxwBnS3OETxW4J2SVDHwzf7OO7PFv5DkHkLFP6
WvBwrpoWIvPK2QvgFp1ezJAtFxyarrb6R15rfxp5zbRNwUVH9LN9FNCSM5T9DRdw
N1YA7TURfnX8WPpU0mRmBSV+7QfuoJR17doTuMJdDK2by1TO4yrv5tNQbf9YFVeW
nj/ljTVefsSG/V/roZk4LsHVPZ3AbOSuYyaUZPF82m6konGA8iw4AmcDXvGWi0/d
ICPVlitfNjDUeGqJFuHrQ1QKb0ywwZCFucn6DDuMMGHRmlJRUjYYE+MC22uVIi0+
QE+2QyWOF2PQ8oyA5eJxW7t6MgIoThrdWyuHEszO93v6B55sco7KfKqlD9A5tQyD
Tmsu/ptlJdsZKKDJKujJLJR4Y9tv9EUZnSkQgwT/iFZ+dFC/jw++V9P4U3rItp7a
CzMneUUAPlkb0+myw1iqggU4cngUV6uYrMCqhSdbfkMKc7IRNBIqnyD7L4O6zavW
saX9KXgIavoSK6LUpOpQIi4kPNYk7D1wTa/OfxcMgJ9UR7yFni5MhfX5W/1+WYVk
KMzgwWVetrjjFUBp9b/E+KP0p5+gycCwi3wyd5+TePMxFhio+ZQf9zMv3WRTYSTo
V2bN8PClIdSw18tzxwb2ByHZ1B/bzvrQPLG/gAvmKz0l0yBpcpw/osNiBs4SGFHs
o+E7I4dOH4QunXndYSfCTk9Djuwlqn8BfgLB+qV4u9/TLdqJXI6AqzUZtLtKtu/w
oAkpXRycHW4RD9iGFKgRhYgCHJazmxeAwqEMPNXcptKZfNsiLMPp5AuhaApNdxxy
y0oudPSFrQyHjH/rzBCDstZdjXCtSNuXDLeGGQKaNVt8AFuabtTRis1tcOh9k+6Z
YjNiHz07RoI80vwwxDbmq830Z9Y+kmxSSgGNu8TLz4gdG8m3ApgQztmk4jGCk0Yx
p7rIyEgkNnIU3qHvdRKvTBhLUWTuTAjYv6VdoTdbrwS2DpU1iXcLFthypfQsLrwQ
vYjA9WG9i+UmvubLjVkW+d0xvtJf5wg1I6YWWm5qWQjeTIAb8vuX9Ifli1eNksnl
wPR0uVQFDTR80pco1Jg9n76itTmHf+mNG5jM0KRLyHTT/prfrTyZtpZKGtf9haJT
DnAPbfPqmy6VjlwPzn2YFcGTCFP54x0hhjRGHoITCoTQVOQLW2NBa2TBqceQuRwV
RzCDzaF2Rs0QYBV4ofpPRudVTHsNz9cIqWy1xVK+r52v1crGV9Bn1/mInwwn6Dmw
gdGITp0e/R33OxKqO6Uge8HtQxV/bhcbcQ9uk4gLM9PtLVaxmLqdpIsy67tAQv1S
f1QpSjDThqRNd4Wt0UIUOgNkNUJ5oyGny/gvFI2DwJHQoKmcr4RzkoS5JYX/wLmp
ljDKzvMdVIJD7zMVccgYq8qhsRvXqLKnEPNszP3dpLOpi6IGSFy1z9s5QCSckRUt
ENb1NMz5iejhrFHMDZkGSKy7EXKcFxpuuDsSLpSBnJmiCFywZR+MRr7gcmPEtOm+
CaMsDAJIXkdn2x6DB9dy2/TKtsZid1uX87nkdbTMTrqpxHGSLRsRczek7bzGkNsB
Kei+vGh4KUpojF//XGxDyyYNwsz3ath7KdfzbOf1nZyXzh8njAieDay5fL4D+J58
k/QWhlgTeFopzO8J/QIspJqDIkAnXShI/TRXFHttx20Y+uyQrg/RHCZA2lCwg5kd
iefGTCBrQSPIcPHNohzTQlV3tD/KR9YlvqQDdhlk0H0enugdidtYiS5bQVqLsp6j
AD1PHv+4c9+nvtvYpCgvsT0ArP2j+4mt8lRKuayqHQrNwMadpnMFnO3QsF6ClYZL
KsS/Vpa1Hg8OLnt9Jxk2M+XtmAufb9MQoXa73HB641/3RYNzBBRswvDjdn1f/0uj
MonkSdvxPg/cMVt7ePCIYvCT/LoQG9FBf7LFvVfoIufx9vNYdJi3FzIkWhZuWpM8
A7lbOp+bTZKbnVj1ybjbZUzoFjv+AAoyFPPr6uALQNG+NQeS7oAEbWspHAfkQ9OW
R0gJ31xKZW+HDb7tH+BL0noKumg1IjRKrAz8m80HUz+HNodWGNctbzboxZ+L9pp1
XI1i1R8M5JIZm5wAhexFYR6RMLO7TiT5ELsEcaMpn7RbYFx6juRW5M4VinSWfjZZ
ZFHaGuSB8GMHWxfEo/w2ZGYoL5zXjur18eOCJGr6Xa/kti6561JVdhCui0i7uOXp
uLRXzooqIRswur8+Uzt45ZxyEKGTFWP/8VPtz68zB7cpWee08zpJwXmMoCalTNuk
XE9uhRBzSo9XR+8Xu8rFZkrB1mlj2EN45mplX16NaRkqsUibb9oea7t42BTNSXPa
h/3T5+0w+afYC2aKxUp+Zp9mSpCGJVWc/iOF0eyLRsmCgmSq2s8mWo7vRvU5MTsD
0XpV0ttW2AarpGowO0w60DG3b5soSfW5Dw7eAnr1SHtN+k+fHMzI5UBBIt9y9Y3l
xbyfh2ZnybJBfmYHPII4CzVY/Zsx6AiUQWFsSwvf2cgs1PgZzrqkg4Tjm3UxiIQ2
dQFH3il8JcWRph+SGVo24REiKph53WSzn+wJGZxoCFnv1E0H6f3kktAL0N66LgQB
BZiAy0zPjj3JaNPAMPLbX1PcU+6gter2lJZWyyfa6Jdo1YWUM4WqjkE6h85lhHuF
9WVSOGXSnyu1OvaD2ND7wuDq/asgW8cIMOQp1j+Rsg8Ov7gA2C8Jq37LUHE/e64Z
ScGozqHSxKAwzCf5Pr0gQrKER8knDfy4ZeCYuT6wXVrLaJJF/XslEwDz1UrANuqh
sd/HuftfLYIlAFm9X+Oi6nEhfwaYRoT1ci6hPpBG/Io2d4Oy0rRLvmvkcKEfGZG9
qd/WXLWBKMOm7HE1H/7eUAycH3eKZu3Ut4TjiTcJie1GrzedBoY9gzZpCXCvsytF
UTTsENaOsqOxoXHCETnF0FmhjcwufttfgLMuik4l7KN+eGW26+5v+ru+DYRbX9kr
RyT+gr1kpptCUsEb33uJibyzVWlaRjfk0DJokn+QHNRssx0CBLHU/qXXngyr++Tg
8r7Rh1f6Q02FFnAEn6UiO4eWxTWhL9u3uArg5cMJLEkxzN4ALxM5KKxLsikM8Z0b
yG7Ko+shSJYU7Cw4nK4QRaq0SA6IGyqQan/HGTB1zGa9p1B1rfL9Hk25nwH4vmLS
ainHZ4DV3+YFJu0zWxW+OmmVpeoLkAPy78Fd8aN7cvRUNer4T3rhiNcWK6B2L7nM
Tj3ctlm9xYyMvzh5PS9pg6341KixsXzxYqKF/OgJ/Jbm2L9GgD60DMVzbquW8b5y
nmb/fRGaaPG1RGgl3dQwdccxbfagmSC3PYZgLrzrHjeu4APEAIWqWzKBwdQVzDlx
K3TEKRY2wdcx+KNG8Rra8Wgkl6PgOuU9nLnYH3uz05N6/j3NO/l81ZqbT3bXpWbG
ZOk9fzZaqiz1FBigV3TeyMlKb8U9GvSaRWoHkS+JMzwwFyF2uRS9kUAaPUWmSk4z
Absv0A113bHboBi75YPlMwz42F/tTNG/+mT9pISAtKfNIWXXCzx9by9nwG9wC9/k
AUfT7fXLoQhFxDxrH87rcY1/XEfZhxGMYBWVJJSmt3B03W+h2jf6G3RFA5iPOVmy
gQ2g52E9nN/vcWAzKsym56FJjW7xr4BktaQ7pJDUD5wXFsgMYSLtdsXsAydL6kXp
eHuI4wFas0SK1JAIZdvm+WiohMZaORhu6GrbUJa9smwCZIUF8w/Jdebk92KTLfHr
2Z0dc5UL/BV6Fes366YUGLZDrDPmvH+3uGE3JUhmlUQLM2GNd+oD0y5pefNapmNI
UOPJzTEKTZ8rqN86D8HqJKWrUSao+7elJ8JbnLytPLHKoS2udqKbB5KMuGv57r68
OHUgLRVon6p3pCgrqYLpR7HX8C2HWKEl1+TGOsXy58JQXmKIjsC3CvE4iTeyBU3g
f66Zd39Hv0R1Z9UCxqGl2CNQkGNkY7jnMI/MCFWY+hzF8D9/lINQf3ZEQETpOxg8
WZOa/UKEE/6JWBgi1r5BXW87zOAQz7tHn6UaKN8ZXvncs6SJyeLxbprhAVre6bFJ
IZi2/aEjBEtpgm9bZrBEQPBf01rY88sEAxG93ZEdEywwMcLw1N+0qiH93iW3ftNf
gfTZkInB06v7oWHGHsfmgIE2rudxD6Fkf162JWLNQg1om8NrFgORovggHw8O9G7q
RiYWIZmOzjx67N67AbDq/7FrRAQCFOp579uiwYoAU9Yow8IJK+EUXGc2u3i2JPlD
iz4l33ziMWKAsEMHYsxrDqJbOE/chHXzDadYpUG45dBC56OircbM+zzmRP9csRin
wt7lki3kBaqYCw+tawyh6DSJEJnqJrIMerQOnBZJljkRuUHy2s6tbrJow43wURRr
4aRfnbqZvzETYXAiYbhuB7ZstA/HxwnBjGnwTi6QvTHlXogJQ+l4pZjo+lzVxNY9
2+/ynkTwSZmBcJCCGK9uM8hM2IeMyBHpjhwUEcXXRDLWwjmesptHaODo6v6OY7B2
cjzcyYqRWUFVyxnnbQHzw60Ac/1zWIZNDF2P8NsN+l/wWX9uTFUfRXvyQJc8ZOrw
FKvf/7EijvPrQ2XMfuOkiutZhpdK1qy5GEoAzIrZ8MfF2sBSljBq1bNc84Qoh8fK
o2cunpQQ1MqgMcojsMb/ws9T0fUcX0lKQ4h5bDDHK68nCtLgdgHOoLb/og+ZZdh9
/gEQlW3TqHS/pWVwfKo8yTNBGJsywYPPbLW/Elrn10LLH36FusfiEQgD14M3M47H
eXrIDBnOIB4IARK79gVvoi7ydqDl4GqlKYHK9LFKlUzHdjK8xwrE/djb77l/AP9b
6NacOG2GCexNgeUblylFYJ9pnKinQ0AEVCGme89Ltv06xDXJ0rYgmkzMCr5c6Jp3
NDT94nI7pH5LYBy2Ljm+ypDvap5zs/uAH4fzbV96NmjZDjsgZbKFFvqiwFRe9u2x
XonfUHrQH4Ett6oFY26HSxZSSN7gUcHT4+xMY0sC9xT58w4HnJA18FUjuno/TEog
orFuCLAgcBtmXciKVgU6hdVcPqUvqFlBoWdYXi1Haktel3YiG6M7YvtE9r8pv/WP
0G9V2N6kIl8HS9CQnMNSerhiGBgciu5BrybG2IF6NrpTTEpy634OCHjLOignsCLr
6d196UPM8rhn8x//rBOrms11ZSTsQ6AQ+Jrz6I8vw2h5vogD9V65BnLqM+3UUji8
7IFzz96LfhZg6FYVL41B3hOLXNY9AO9X29b98NaulGw=
`protect END_PROTECTED
