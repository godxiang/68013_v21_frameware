`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+mHWMVvCbMh+chJ/G2qI4FgsPdbRNnVEjQT5Ub+gmLoPVU2YxPdVp2+MO5ooyw4
GZEBQwHzQ2/8UlyC3a9cjLF5gDUQOMieR1mUFDpdUSSk+jE5HhRCeo0zWw+qBh/P
p63dNHhxuTsyO5E9UAyFW5jcV7SVSWxDvFk2kt2wXc4zVz5bvJDzn5rCf12SkU4W
2HZGVVVBFFpCuZ73QGXOUx2Rrg7HEVnfEUuSoLez6+cKgHdq3jZ0ozpuyfEKAEE9
ckPzx5fFI8QKzPB7S4+XkxhFoTqhFWtb83KFzprROAV7P2laUT2TejUmpYIJn59t
eCmdGd8m6dYjSRxFqHBcAgfuZ2M/GdJYBdXEDNrfR51TK8yYUkKcoOJ8QhFqt79M
wD2i/xCNOA87iob2fiD1EJIHRmBWrgl7fyGaswsOYfaL49DWtv51r2CflmuIao8x
2TEg8qRXD9VSZWsBYd6Lbe9TN7n0TmNmJWZf97ZRuVEAvkj0Vwy2l1jLIJL9XRBZ
N4XlCYCs9plpR2Al/CL/Q/Kro6ni2D2J/cxgQTyUmAgTkX+mx5128Bqe+UMI7uEn
ZbK5Uo+lYuyRDC7eDLag6l/DWAHX0ZIjUurU4L5mwcldhkZVIRlFaIXFNgrExvxR
HxNLXSN4G3TUwfFxfT2nzEGFj0tE8KoLNfrK8Q195c1AQi48/Br7wbhfCTv1DD4w
x3i5nzVaF+VZjMz7ZtKJ4h0XGHUzVY9QQMxGJoe2GoVWw4r4ePTPavrMKJwzeIbN
jX74qfEd29Y9NXXkMg5c4EWmpqs6Fe5COoE9j5vn/NMc8+mHS4GuX9aiPWBk0Vds
sgTOaLgDqCKc878FTxZSFrGhIyOe2KE4+2HR+syH/OR/zkMOlqKCpUP4+LYdLyO7
1RWqdS6p+MkeWscTzSCHKUnQrBWR+kvIzc5ijSJjv3PRFk3W1QdaFxm7vm9JLhlH
lKYMc9O8+BjOfDkDZ6VmfR7kMIS2+MxBAqnQwOV/Id4m+x0ZuLUbv8CFVS229XQz
rofr+zDlG1pt3DSiactuiVn4mklz4dcKBJkFyleO4iaV8bYgga6x0kzuB+BvObwP
8xV+Yy8PGNkCTaaQoEXbOXzlzLzmHuDQzlf/IxoV960QaWnAXyObCs2cEUYXIqtc
wr5xT8RGy83KUpPH1+ZJj81r0OPjV2ZlKVQmVcPB22C/glnOybVhaV46GOCtpC+O
TTMCDvpm4ex5quheicw1RlYCdh2dOSGrSc06ddRrqAiA/KN73IHp41lT8DHfkxN4
gy7GOiP+I/7M4VV3624+RgINvFxe67w7ckyLkvJkumXEHINITZAmbh6ahnlpzdlw
KZWuSIFqd+t0UKmz1ZXdM+Bd4hDB6/ppbOyegEoZzNFwysLsvyBb9HbkfEdmNo/b
22raRczajjAz9T/+ixiJULGc5fk15pQWrXdzFoX8aY6Mn7shWjbpuFut+vadushQ
gpqNteG1MLgtT2Ej6rg23R/hZd9v/+/aPO8Y8e7pjVpyzuOGhLo0VHj8sLt3MSNk
puffVKwG3ECxDk/4lb/4is6Nbypmeu+ExfWT7r1XPvIzgpQCessoVO+afL1ex9ft
5Xk2XKaTwD0hTQdI5AAnjpATDsSQW0LbgkDrjoJuPoJ6z3tcLp1QqRR3ssY6ip1b
3QHBjSZL4sgsl0Oo23LtwzO55m4+h/5FQnQy+hsvmBVHX9V2c1Po6SZoZIly0+lD
LXpdhJl/5hfts7EHDemLiS85owRPqk8p4n5ZFcxShKXsu7kWaXkeK0XiEDZIl3C8
lss7naJF51Qamm6bLQim7SAkjS06FXX8tQuYKEJcXW6B5Bfi9lcQNU/WIdGnpuhQ
+aiIcqmQMaWqzVr7t7+PRn1hEY8sN3MYa2b8ShHSDS0d591aB1uGRNaRHpS4LVz2
vMhQYuZVx4+pzwgpKYvYAL7mc0Eg9xdHhdtwLjvhwjo5YHlSeQd9LgovBRj1cAhI
0Ti7/41nS8BcfHb1Nxd2MfDpfq6otw7kyEgeP3Q+XfveFFzht1C7u/niuInPDWiG
r2XLuFx4zPncVBS35qiSwDrwc/zOkTe3CbKNUxQGxPfx2Dt/gsvfOyGRsOE1ERyu
UfRwwzIoQb9WNSYDw7dhgBMGQBFUnoi1HxjnLRcJd330bW1jmx4viFdQrhAhp0/+
SA23BlgIXDfgjG9ywBPJrukVgIM/R21KU1wVYuiaNgSnrNFYu4Xpq855lecXNEvn
CxWf7Fhi0qzrHSCMMlbbsHFHDaJjBk7oGkxgmhyqpXaxXDWxRv84HNxyq33oYfH0
WGcEBAhh5DzjK58NgBcAv9+/g/BZ3u4lsni6IIIzm5F2g3NJgupPmNMybL2ksHoD
aA4SXOOqbHZZWmBmNtMes93b3k7xn4LIXWZfQSc5nXk+oN1DGfDe9P8ohmRitXse
EJEaYJcyyUwP3oLHU6Bjec8CSJnjQugdlchhrBV6ABBkQf6J69XERdiIwuYZsRLG
bndkR1cv1AUa1aF/Ye0czSf3I8ulayfoQK/KVy9Ec83Pvt1IGsEhzJyq9nltSSXu
+uzdvE0ISS5IUIX2eQC3NrxQUAyvXXoEDUIhwLpXZYbw1ZrrKPUM5zNDT4vNgX92
HHLNDTopKSGZkH4MOVtBWgxdS2M7IqhPyBkrIbazkejAmvkEO+dUG1p8GaEIUqKQ
7XPzdIh3VE4UWWaNdOdEo57SArhoNPTYYPdyOLghSwo+pHGPn1hmAiCL9ms/taXK
5/tLA3OivXb/PZ5A7ycoyeG8bwIKRDaPgkr0hRwRjTMo9CLPYkqLunoTRS65Gu8h
upO7b3ZoBqHw46ow+WrKiiCEl8uktbQfKJMS3bLqUk1KX+Z6AlyOENDwEIAViL12
1QZtgFIwbSwAxiFmM28SmtrMco9qiB4PeppHJ/2PNLf58MMcbb5R94zHK2fkt/Vn
WLlGp9+YKRXQ8lCxNivE8NwxLnEu6+/Rny/bPIsxFaBn9oPLkOQ9M9Wv5xfCgBb1
d+z8HJxOhrifTtXZX0akrz+BcEtEdVJi52/uqmWdTyR9VWYjjYocsIzBfIc/3s2w
loEF7x39J/A1nbpLQgM3eI58CFk9xvqkm1wjqpMV67xk9FZEgypdKuXlfiP346xX
3eZQVLdTBPUZ/tQdLv74Xg6LQJc4m9LZ9g4BaEbkvn28kMexwCnSzEbkPXtQs0OU
4QVQTolmbC2HXlz3JqaLJHLJAHx9sTZjWGYP7cBQU9zuiUdtpnrmVFlb4a0TknKt
di1PfN543C8HdhgB+DC4yiCs+SeqFvFNkG7qCyqpX5/Yp0/AA/pP863GKkG0T9tT
uabcp/CX85P/JDqi9kNxsuVxoV0hHnCGg8a3DCbcxBV/RSLjUshV78lGmFKVfeVl
in5aZlpveuCmidAde8tURRinC/XvNCJ9Ja6y02qBFZm6y0Z9D5VhNNAXmSYdxbkA
1b2x8i/VFxtQFYaX90/+Nc1YWUmn148kpw2dJfQ0p+QYg5pVo7K63WNOoepdKFBp
whTXp8Jd0hAPtHLPvplb5kFKp9L5NuPziq/3NxsYU+2lJlhnvnB+Rsj+yNa+knBn
aAqDvZuVhZVb9yxi1YttB9qZTnrg+DySGyOX+1WKF1z/CDe8aA3pjdAkxrZ3/eX4
xtJaPJXEouBX9q7InwfojPUh1Lrl2DmwxucwWZ7HdwUC/ajJ+NHYar3h353yAcKn
e/g9u5N6spQ2Ww1R6UAj5qi+6t+91ackMDR9jayJtwyrHjPNWRsrR546KHyv8QHr
V3i6l7UFER1ZPJidOH+7T1qKZwm6rqzv8XY6a39euDuKA0VM9KgiKZy0IY/u88Ky
Altb6RMjAwOcmRA8Hyyj62QFDuj+2Hhq8mrTxbHZeHNSc8vpqFAf9EAThy4lpgjo
+Fl1nXSKtom9rd0MD4iHoJSQ/PG3/M6bCC/7LKoRhGDRWD9bYOznsxCmI8pJ4y3N
ISkqH8ySi8HPar0ZRgXnu5DRIBD6W5sTS7Va69nGc6raNjo+ocQflyH9n2zeCqpL
yvf3W6BWcmuVDxsqkZ+KDZCvXA2+7iyy5NBnTm3wxLz6g4TAzWyo9+BkmbMzJFpt
+2oRSFHC05HTIM9nDeGDwKkjawKvTFCmekRP8d/NVOg74wnQaK+a2vSgV/HgewDe
F3iCbdBEFfE/gwabUqPJ7XGZTFXI7PgTGBU+ec15Uw9C6ZNg+faHOo55L51RAtrj
xI8Pp8Md4hxVGoOr8BSt5TdIHu11amVOvXGoMiGB0QKILprvAR6FTy0nN85At/Ob
QXxvYQwGz0pOMIouAsFaJO10VCWMS968PCql8x75YJI7QK57MVLDyzN/1AlrBnSk
5UxI+ES3stGJeu11SOz3WhWzGcsYyU2wP5/PhFm88bxhsd786VYXy6tvWcOO5QEE
UfJ2sTBr6w1vehmpLwoI+FBo/8le6TptvgwRdz6yCeLpMkAXE4TAEa8jRamFxaMT
r6sNQBradzxB/1en9wFqvZEDHQDCOb7LUVfp7wst66qvE456yHUjHnP9Vii4vDtY
ta0/d2uqHD8isaI9Xhab09sqFDUZV+k0O2i28p1dKqaDb4Qsk9mwB5pVW6enca4a
/kZC4Jjxkc8ksdJcb8T6cj5N8YfrSeYFoy93CLgz4wZlCb0edvT6rKntgpgOJ2Gq
vi2XDdquj7h2rrI7YJC5DGOLaVaZveQSQMD+n2bSQn71bEjBhvhe/oY71WhUqXZR
r1YmrZNPfijS1b9PTpQmoqxDz+a05pLtnGBSVF84MfpOfKRzto1psGx9SzPJKBC2
5d+thiciGK3ijUkZtIoSeiV58WMvS3yWjU9DsnaZYHXwMKrbRwN+hRKLmKY0V0aM
G40KTgEmQXNLECQO82lVEg64J9RLj95BipjDQn4JpYmjAH9FXzmwuCf45VvGVceo
Y75TSovWrbyBw8SXEc8cXX3jOxhT6boI8sUBu0hp2nL20yc8GczdYoPzbCJ22G1u
Bp8e6GQe6QHZPgCQx28kQwWqXxyQnd+P+K61gqCTbFVJ2LSW/tLbWEk5maZf3XWY
hidroVTJ87yuoO7Uu0GVI1X+JC1LgevnJQd8FpX7vw7NK18rXYvdLkwNAg0F1B+/
cczKiAi5Iy5QZNcFDVLbmdaBL/C5EmrqzfBag76+4cv9SdvThhnf+OTEZKBA9KS3
xlpq5hBabnC4LALQEQtndfltMPQZvUrJeh/Rnl/7cirE9WuT+ZNPKsKeQOKka8ZM
Un/mrWrkaUm3tHiwOAI5IGR5A81cjiconwaojkCRVkt1366BEXeY3UeNHYGG4v+Y
lEsXFhsfCmWa4Yd5qvHqCeB0msnOBP8Hr/A0lTw27wSE7+dtUiynLHh80uaVpPLj
u+TrR/1Oc8LIP+mH2BdAMzEgcQrJKEy/0oETWuZIJltuGuUWQly/fJrpdvH2Vq2s
RNlo1NALOEHOV+9vMAsWdo0gpyzKE754MaX7afpknKIK400jjD610RpJFZPuClzf
/572TdkxcIcfqyMCTC5kyAtQbikLY1GLN1+3XTdWbTMe/PxPdHAXTVCL8XJZwNFj
tDoI0CK+2LPZ12jrEX3quRSdiGfXQc10jRFoOUHHMzoAlwmyBulorVThoBS8Ll9G
hzhyLHfS8psy/7PskM3xQAKCx5OYPvQGXKPx2zRtC16S6RjGyLPQDRygPKoUPOH6
SzUhL1x0LDZPRHq/B67k8q/2NeRF4DF424MXZRTNiWjB7OjqI2az1QiXHpnv6R97
A6+1zG+cRauRjWXzYek30jWp191cmihbKLtPmc6NG1gjy1puH01akZbLxLrYXvKy
HXvyZbNpAz9ihrQk5ezmRFOabwcspXnQM1gC9TDC9Hci/QAcHv1rkuX8F6izHkPB
/EtuanvJcp9mhGkK0cx2tL94ASyovhtGFWPiViyaBP0CYP6RETRLwnUbXSaohCdS
W99DztM9GMYMBtzrF59MPVys2muDIcKvd4+sxmQZ37VHhsbVuc2RoORX8nAK++hZ
/3kQnDJR1Gj6a6abkHSU/ikqzK0/hEqwlKtiywzwhdNiu0N/xnqN/BVbCrTL2Y6T
GAVM4XbWS0ltaaeizBVRdG1fvCDlKxVlBJJWShFCFrvkVAqwERq5ij4oTlQOOTI2
j8Eon6fCM8mmzgsjhc936H363ShAN0Tn0UpynMvYR7lMlQ3DLRU4/Bq8CTCcAR4J
0J5rJtqQcvBA2AHCaKutGrXz8nPufUYuFQ4aEpCG0GCXlqICf81jFawY0o9RKlzH
XJ7BTKgf6W5SBCVdrl/3kf6KLl6HNs2YrkCjR9RseooDEV8Y/VhsXGZSOcPRWXSe
H/H9ngjgCVQmzHJ+MjGaBA3pHcxI9Bpt48u+AjDVIMRDrU/bM+ZjuGu2NyTt9WH2
RlNRJw3/msYi2mksLiuEAb7cj6uSn9MOJkJfTYJZ5bdtVQ/Ufxta8R65vflqUTFk
Eq/vVZpQIeHylEtNIjDWgbrWZaxDRPs2PAL7ugFfOrXWGBl+3tdGRtIrVMLpNEXI
hqLqBqeinT6X/mbSrmTchr4u/Y5F3x/sD6ZWdvVV5Bexfjv8KLC9Knhn3P8d3IYj
6n6hZIQ24LVAzBbKBD56SBeeYdK5R/47qpyAbHdvXoqkZDB9dbeRRR3aKw5RPgK8
gk79UpszDXSWTjZGuj824cgbRC1ro9O0eq9DzyIO64CKzxD9r6cKDK+mzyDA/F0o
3JG6j5aMBVKJXiJ/Ke9mMrJDZdbIigEREypCvLOzwffYaM2JgSBygO9Ft/7gvAiJ
nA9YDNMLIBLT3EM+rC48NW1rgEhYtee+IOFzSe8UvfVuOpXMhDJ+Q7tW9zbfOT2R
B8Zzv9u8rQx67Js+0I5nupURxX4bf9ffXHb927wGv5QqJU4YN4MHyEuYELD58Xas
5zEjTY9604TYjpf164BUA5PaNaDOq4+F+aIHZ8Z1NvEwOdXgur5vsl8kOJwGR13D
Uecy5bPEWq8m6Lg1GqTSLZNUBpq4O5RO4Y8xn1AtmUeIjyD++4931n/v+jjVFYhg
fJLOgIEwMLH4MKSRhxBh+/CML4nde6kcpT0lmmvhYzmqGQS/baJP38hivGMTWNdB
KtkHiDE6f3ehm0aDpePluOQmEuazbjIN0W2SUoJWOchwgFgRv+FpgCsR6IJG1wto
ZZrOfXwG7izq66lcnAgLm/4WzLYaUMnrfZyB9a2h71oQwNiY6bFl2aNgD8kJEri0
LLC79TtUE0d53NmWY1PT+2vRA7GnufeQQ/vNm1ineAp+vWNnHQUe0Bb+WrDnk4AP
ga+gN/Bu3BWa13VEmDTv7dc61qEVrMIOGtx79wVQS1y3vKWVo9OwWNo6VQMLtGbB
JJZJJQTWmmm8BSrCJGL07PV9L9EId6zuG50czT4hqb23vRLmk3dEueRGup6cMAlR
UGfURI6gddjk065oiO/NY6OcTqZxKRb/zV3KcQVR9cCr9oVbIctrE3c4FY4fYIkE
26lOcLMbQ23l8VAezKL5+i8KsW1CLQ6Xp5vC6PKb00S0hYUQLGxJ0jazFORG/HA9
vbG4kYM/Q31O1vNt9z7I+xYmN/ZpLrFPmitzrhlj432BYL5LQCJh/LgoJBTr1AUf
n357sguNkQ7cdAETu1KOXHITRLpiBaK/qhALt+yfH8BAGTjeMANWD1hoVlSM+AD4
2ZtugHJkjnau+PN+G/iYXv/kFK+jFaGBrLjJxg4Mqz8esZOQZ75NsG7keLAqyVcW
FvQqKiTWs2sylEfr5mOQX+Zqe0pq6QD/zLvm42KJEYilylnE5CX0aTmf6v7UVzY9
0jEKZYCjzcGfFsRfTLe2z/DTihrcuk3mlWwicOpygfwBFo6m2x3L/qtu8pz2I69+
zKQNLLRLG0ECbbVfSDZqYVoUOyyR7InfU7IxQpHfLsjguCP0BNdMgqx100F9lAQz
lZwVcWCeJLqMv7bgF39FVRvWB+u8rq6H548N/j1wF2kLksqHl0GjqqszgtOrW7bI
/zIg75/UVLChO7VN58kjGRLxZ1MLQg5Qfb8/uEs4xk9JIbjkS4bUYUf/2+OZNnmQ
zy7LEdTkyBk9J9OfJNurYTI2PiftriDbLEGVknE3f7767NhWlu80keMKi1PJElYs
`protect END_PROTECTED
