`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I4DQ8mghWx5zGuwFOc8aYrU+srKu/7x+Sngxs8+VzdhgOJ6fVLhiDe+Ouhdzoyy5
4ZXjQmkoUFW6EH4xFWXoJxr+NLnJvEtw8JxZ2/kMlrdw+0pFA46nwBT0bUhvan1p
DsjtEz0bR/L3TIO7dG9pot/1ddYKLg+iMD1fhtLvO9oZ8hrfwTVFsEt6WFlYFJqD
+sWZmWe5/Sqy1lPuwjd2u4wSjcSvVnClpZiLtYPgzLuerKY9vD0/lW7QdEEKMP7B
wYA8DaKwcmrH5QHbqni/AqIwGGnL0vk0O2pr9/7KCdkaoVC+m8D8XG1QFKl5pOaD
5Hw92+ORJUGFnh45JoZplQWvU8hIzY5v711koY8uuI9pDpuTYl3VAySOYw96pvqs
bBgXlyrNhh14nZaTiwGFD8R7IiQLaMvACWT+1nkwepCgDzwvpSQZDrJLYuLijozG
+zeeioMBsFVtwIM6IXY/lDjRNay4fFoBSVA71ml2AFhzAlEwYIr1qKuwkEeAbn8w
OWnac+9jiRgmurth+yDIga27qs0gexSN1ZGHfaJSg9oZDt/XnaZXFy+tXfyrRWFD
iHjcQglsM3UADKll4PKE5TcMC1+U7l197y5MrPbH2QFHV1AG20Fi8ESn9MHhfJWr
abLQPNO0kNE9WixaD+VJZvE2glXmwfEo0ht0/GgSj4+Rv0puY13rSBxHmI2zrR/5
7V6gULRbOuX3F+3Zb+nT9ctvd+WtnnUYZOWP9CjtaZpQ1/Hro+cX//sPu99HFj4G
dcqzG8qy4t1umhVJMkYGa22Brm4wxnVw0wKQKGE4vO5+a5zzOD1yPvGK6WgDxFJM
mQ3oPm7cZBPZ3RfJGIkCJMDGkycpXLHNHEg2y1M22shidD3IcyKbMnBQNX/DBCoD
YuoZrqPntFr+caw+NewOdU8rYXD9QxUOqBOKvE93dG7UuLVzLeJJm9k9JaQZZxpC
bfnNaz38HgJyXje2j4zZjrzMFtLRTpZMUC57V2TPvyOim0srbswMrqwaMMxjANI6
z8m5IdDj9mo2HEVzYZlEeX2ZbaVNKe+B+NDkGqvPT+fDuVHpVt8dmcjduZa/jVg4
WWvHPvQ+qCSgxAje9TmZsnvhxhysxgMseaVlmwK3b5xFx45iSsxEkI3DlE98xb/4
eO3wgZ7VD9W44iI4b+rOrMZ1s9nEjyMF0tk7N6MUb5aNMkXvZAStk0toY8DnAqO8
PR9S89bmGYzmFk7hKKNLMi5XahHlQKLYn82Kf808zlGaXZaD5uL6WG75xeOfnjd8
h8b48Mhyt7HxtZX0LcJo/PW/LvcEJMI+htHkkLOSEdNhrZovQ0RpjizdXhOa4WYX
yjQmiktySdYRr/vDHIadDfKzKCvTppla/FpfgbNJ32NZAmGiOewqxKmeJUOm3sLb
LiF6NMyVWtHPYALs4kjuBbkGFBBwIIFC5GF1YVc576BPK9gi9XWCmwnPkF0QSz8E
gVwzTQbwHd75lCUZ0Yr/9sbZWS+wQcZKg4CkJnRmGF32bf94RD58Axjd5J5yZatu
JqKkglTO8DmVUukbo1BhA8/ehjkxjHBU4OF5gst+F/2BlQ/hXa/FxhFHK4oePhr2
MnBo6fzBit3GtfOaDwb+qT2CmtOPNk2iph2iivgtu+cjhRQbyXJbdRKqPGvT0gaU
MpPSLpMZ8pbDc9YioQS5u8iOIQXNG/r8uNm39K1r5/LfXlabfI5Z6xYgPv52eWGH
Zz6f5bsZ22JsOw48OCxIlmDi+3WaG1ZFDNrJtMNaZo4ZAGom4Pw4DUQBXybQDheb
OzGKAITV3ktp9k1SZKphrsCW+J9lXcL70iLd0zSh2ALZdFbkWCLl+WHEcw6XOtz7
UebLhvrUCr44uxQFQEvTuk3KK1K5XTnn2L5xjDvKqgGe6/36sWU1/QRhzsHXUUPE
VEm6cVNcEajCWV6LaW51aNiAuRqxQpc76XvtnsNKSRF4ypdZ14Yww3nAAhe4PYPg
Hi/20fbxNgNFxUmPar7CkvyKWDH7qNYlgYuBNhmsaIqIqc+HmLlCr8vNeL9u+wQv
nRRt9zaKs5FDtsuUDuE4Vj3shajRcETgDCZqpmyRze6Q9V4u/JavoqGzbYfq2GMu
ZzCrtWImqA88332cOKUVwsuwgudMvv1XrN1Oaysx/1TeLpT2UckOXI5HH5u7nRXO
/Jc/Zpw+LGUhjF38fUPE9DeTMomKwZqNRCViK9Km7AAoOS6HYGq93WE2q96FKS3Y
8gT2y9zhLZdH8ecfzb31W1OqCFRweK/IakflbXMeXzqcvLDHPAtbYYbG5iQjQR08
Ti8WemckJNNhA1z0NUpOrZEmBbUL6duW7w68JJwx/7XU8fO0Dc6cRBaPj8XvRWmC
dzeoBgI2wyaBz+NHqSKZvzpN6xvGCb+J6UPHXB6oCPVKL0rvOvI8vod5fSnRol4j
kmAIGmQe25nlOmUxVDTo3vRGqcWoHQujtQjmhsWg4Xwen03Uc+W239W5CaAUzJ+N
/R9jRDTl2RL6QVdIDCMBR6ea36w4E2fPEcq5qRDY2w0rRaMPs1WvhiivflPg5j1N
eiSKsLYNOSuZgfuLqj3O/T6ZBh1BaAPAz0ZonA3iSisYfkWrRQpCXlbtxWT01wrA
PodM2zNk0rRZdspyfHbxagz82INad0VXcfjrJBzXnDKVtD+jfp3GVzk7cbFITa0S
vEAVIYO4K2MjrW1H5Jq8t2rWHYym+p1By23OGdsNEhq9WMJoTAKDKcrcRooLksPJ
XC19NUNBGYr2rvMsb6L8ifziFw1mhS0uPu89JExCljvegPx48kLUw8sEQIHaaX5l
HIXuEc5youOCWu7n7cOnBRkoHBSLkJ2LhxPMRMzApxWxHHqk/ZmNhcGnElQpkQdV
9pv4B6+TPige/UpIZCFA3WUSB/fY2hN2kA18xt9zdpyyyXib+ll3bgcDpcTtdZ8L
9RulCykMReixonAHqGUJHIWuCvrFPBNQqiCUvp7/7AEyL/0vnFS6ZSo5lWbrIuiA
C+RvZTMVTsLnyNqmGAaiyh7qy30T7Ua9Gw/C+9Za0TbTH3ZTP+o4VZByRQJ0NgcC
1UBC8ZaFbdjbBrJJ/pPpm1VxKPpPJvjwME7X0xfmAimIPpT0+eb3BRIvtZjjA6jk
BU2tPCciFH0SJp9nKfVEk9BPCLUuWNqEdXoK208HP4tcJ2I7QgAXA1rt/CuM6FGS
5Q9ynnLAwdqazSzIzoR3jVmGrtjDMWmFnhboh4sN5Kcuo/Bg24JuCIj4RW8kNAqN
mnwDhTmiJvQAXEMFfcCK7YUqFIL9nkN7AQQxy+RpOjzqbEbiaL/MKD24NO6kF8yv
u6rH5+BXK/3CoaebVIIEfmUe+/Rh0UZhAL3cP2WLH7vrRiI2PsKjqFivqXUzsjWz
KqjlNiv4UmBNbr91+XPHGeopsUfXsJO4tLbstzuMmxSoDAr4w0tEf8urFmoIitHv
qoDbngPcLio5dqG/KHsU73pVNBpLeVq3WQyhs45j0xGp3lr+ZZ+G4R9nNT5Yb6Q6
4ntYpA1+en0+MAstoLNL9mTH+Kqps9GWSHDwyCDedvAIq3QSWuND2C+5lRa/gmiB
jWfJkSgmiKoES/8re3V36tGxRegTPpQYcgwJsSMUgjR5PlPiwrSqBN8rUbubl2G0
wdAZFEJNj9HVas8LU3JWtuo6XD7jg/6Y0xu0f5IHWm2d8z7v5cg6uGJUQz0P61LY
J/Am37m+dslo07CAmtasu7jKVUvcj+MKNA4QL0mA2tW5mJ7D4O+wzeNh2SkLmYm6
6sO0EOMJuVsq6qO8bq8kimCaoIo48UleRR4j+wCfME3fIrAE7Sk+snCPQK9HDdyO
+a212bEpr2Zl/yolwZDG5UaaXZIbk3Dyt6s3EyrnM9nu3MP0l7N6qInewvbYgiaE
bqf9SQ9LNAwmow+7lK4eJdTGepp/uIdrMqD9M5NS7ikoaRXYDNyc80jhty82mVhD
H4vrn9u/R8w7IbcF9IwXa47Yx3QHvUMsZfiogDGOi/Bd2bw9jVohmgkK4KwiuN9x
GDHGzzrze/hpO22dh1pK2/kFQPTrhFu8Z3RLePMXcoNRkVvnTFg1567rUe5t91/T
7UKaD6o3GUKRcZludi6J4obkjck//zm4egOPYRTSbU2aeH+6uzGhnRle3jGncf9g
xJqs3wF4sP+MryWrzR91QqCWFXvOnf95PgV2TICDKupI6QSFckHkpgbnkFeDqAZs
62oiEg4VTnK//l19E4UWOUiQv/fAwVI2AFTEWzlaJ1f5x75RDscGlH4De1ZX0B5u
62NUSeOdSJBruqt8HB9MOp2LSGm7keyZfSjVVL9CPalpCfWGceUnFz/PwZyFv0ae
q2j3tBwjei3Us5WfRIGjdw3FtOnI0P+Hp4V4qts8DVJPi8MXYBLKCgcg6zVGL/K+
77cMjyJMUDQNtdRXZ4jB/NuTvwTpQT6INMjjhIntE3krlEo7E+yKmm84Yf5cZev9
fPOO+k2TLiXj6K4Rz+x6INDolTCJ1MkHmSoC1ChnaFOhcbpdu6996uxq2LBGsc2U
b5w/1IpK7GW/5b98/J5MECNN8BJ/RA+xMG1iaxMZp6p/ostZ4RxLvbaFK7jcZgkp
ckhG6ATnPUKIs/1dKdBbn3DXu6+LxQLdjTPGIgkNfZgBkA3Wa7lZtZi6b0RFaTH3
Xl0gQEVRFdXUbHKKfLrWgjbBRiwseJ6mUW0DLGdK51lty13nNgkt8TBHZKlp2bb1
oClu2SkW5QtxdYh7blum9L9GuDhcdmnHvemotSU7GHnWugHwqRezd+ZYRRCEdtXr
QMOEqWNJRIu1PWGG5Z/IE+sj6xIu5tUrP/BRQyC0BvJW8j2XGZIx40hWmgpOYTSQ
M/7RFbYtdbUnjI1YM9LlRutEuMki6N3SYA4RICNxfEnMCtUCDSKxNIlch7CCfPm4
4hBOIQCUYsui9Px5JZGsyFs9RRUM0PdGYM4fR9fpbBcxxt3+BELMn0NteHFxJid1
P27FdCE2X0Zjl+Lu5w9E6quBFyLsYETQMsc8N3Qk0a9iNlm2FLmn+NoyjvN+iRMd
/Lekf7WJGFw8+4w7odl/IuxBhBX1UIVwE6paC1AOyWc34lIjtKCOODZmBpTaCf+3
hk5YlyWJuT4PA8T1u4U2R1r1oU1XvyfgGg5sCu64kPsMK51OuQwdkOtCm22rrthu
MuOMCMXjb/+zABPFUSj30j2XsGyl73jS9CuCN4lXR7moED0NbICEzZT1l0zy5J76
iDI66u/5aGf2nHh/CJufgaGf17h8pLwd9zeN+eVhBLpQU2aODgpzjuaTq8xxDHv6
VHdj5XO7N30AH0V30GwKRnUgKrhSMurlIgfvtVjpjCaDdVi6BwLZz4X3sXzPv/F+
MAYgnjW5QyoyJUGJ7y4saLs1o/WcLlqLayzznU6tGn0+eVMiL/91uI6dCDZASIQN
QQLcejTl7ERNDG1AC8vaMUfVKhRYxALc9VWta7ah6Zd3VRMaFor+HefUtSndcFHC
8uHCv2u6qwIGmhs7D9CWKLuyP6er80gZvc2XzUiv89h6DnLrLmLCheGzuRov+aWY
Y3BaiBteoZ4lItjDOAvU5R4QL777Vd2qVbORI7GptLO9BiK8SORMU41CWmvCFxWF
b/ynBvFnHZptyyFMt+3ipFuf82b6TjFLRBaSESwddqfLWBJE9BJ/pua5yqch7IQ3
AkPOE1+0UVmwIp1KYzYw9chY0K2JejZtp8gpp891xYZ8B8CqwJBA6tSUijjK52K6
zjqCjkYApJzv7YST4q4A9gOlblKe2PuNcwBdk9whR1tV8rbul1zWimJmYOCJ1uqe
h9JSlQsB932/Q5HSJyS1KhW4eH/8paIh7Qz0ih675l79dfbYNrzSOXVAHnDtjX5a
Q8cQCa3qujxxo14NwxC9tWf24Mae8c4Yxsry16gELA2hft/y5yUDfOVG4PaWfb+V
m3lpkevj09yJmLM1OiGVri+ptlzAiIJZsW95bxG0kffQPSUOuBn7u0q8NVwZ8h9j
1w35e8bShc201z3jqivXRGOwOCN6KOru4eVb1wYSJV1UrdT8Oum95oqb/6L+Gljs
WbWV/EnsmMHJ0Nc4Fg0tHkv41LZU+2RW4iUFLmjjm+95emzew141Z7Rnh7fhE03C
zqPM86aiiRPHpEfIgej26zkcGvEzSnrYYLPv+u2GpQpnlFXRA7heTBcYzo41jRSq
GvmUMjy+3KxESFWbJ/nDZSbZwzDPg0knsJKwoez+gg46C76iPV6LofVcIItDfBwW
qPEHIjiwgbFukJJ/roxLyypKuUxTZ4ujz9NKhxRjxyKoffkGMGIOPHScNPQq+2+H
2tt+RSOfoIbd9Yo03DE19XrKlmY5F3eTSzOR23towmvVx4t24u8pmwyauWSJ/HBD
zQZBwgBR8++jSS710K6psIjqU9hMEq+dk97lqMKyDcX6s1EeJgV2cdgnRtPh0Otg
lLpZXfTjut4BlLGsPt7pWHRi2TCcBes/Wt3PKGL/JG5+vw25QfGbD2k0YknuSO9h
+13J6H8W42xmwV1wPzckanOpGKvUSNT2nUPMwa6qfXWFLy8LUBB/f1eAWkDoCgoV
TqOVSTrhYn19d+ZBTCymWWb1MjP0mIyN8FY18YwWc90Ex/jYcA1RpsQmAhOfnIm0
9fGzMOydOA8D9NYuW0HhTYKa9Z8nLicrJYm1Q0glN9eXLTtH29+QVl9AWo4RX/qD
ZnipcaNvwvvVcMT50dmvmT2X+IAytu/n/JH+D54I6x9NXVRjciBs6h6YlUkGUWOH
NflFJuhCnWyP/g0FcjlmejMJkMrWY2pzp/HiiX058EKeRrU/Me6bBMXh1xV1c/D3
wATRRau5cRAZYZwvf85G6hZ0AE284qjVmf+lUfzlp/3LdZsrWXqwdFhHpfAjgDmB
4KrtXY7pLnRh/I3awHv1TuAv+1wg92RgeRcIB6VpmghYllxdWbK0peVMNdjCHYcs
ImNPkUe4aF0LwI/mkndm/rXvZOFFhOgmNc+AtU8WUluze6CLaezyQUS4NdTdW22o
a8ln1Hw/46l8mfE3/emsfWK5HaHTeSd4ct6L5BAOui8ATqwww+lP5V/7w5Jl4Bu7
7Ittf1fTxNqsSJZavYe56OHdlRnbZjkndfRLnrL5G8IxCsY1SxZViz05/lmSuAz8
Z+rtNR5AQVkKUSwwl2h8auHUxYf6F5n8zP6NOYbSQz4ZJlTtYkYfwKa1cygOpXeg
533tlcGrZnYcVn4gPDtUwmeND1GDxkCy1phet2snZTdYttBnAxY8W0hTtrOomIuZ
Ktmvk/xkzevUllF56AybfivvvsKGZTiuKnMnRomREOafvIOZ4CkGa1dwxIlEkhuD
sGe5ru1ZRNgEgeUTdvFcSSD89ErMQuEFCUoatov3pwTDWrkkqpjBpjuMzrY6Zb9c
uY91KWFTvhwoszJpxQRX6zr25bigYY+xkW3147eSxp2CJVp+7pf1AnHVFccZv/8t
PAxCpyzVai/KFKtkNCO+KZFwuZ6quhdyezGJdtNLs/t7urgmzySNyqCs+FtlOYAp
vA+cDZSZQRWBqOM+/gx6NH5h4nzMBqVgYNw+bOgsy2n/A9grVaBJi7xpIC4ETkPg
4+eoo8ijl82MECCtx0e8F6WOnW3ExU+zkq4eqO0q9db8pI6usJvpsyc7/siZrt3b
TZ99OiQImQKOKUcgeA8YonoZYxNYsxJ73O73QYZJzS77DqBIMbnJJfRRs6L9fTQW
e4YQRFFmRHM3We58G/0WPTExdQR7jHtVXEaYH8o+Ez3AvvfWtLLeRWSNfuTd6CzA
s2d2pEophZ2xreKHp7yPncKOirhitDwHd+eI/T05P6BD38hdoI/N/o/Lv0CxDcGV
gOqVXnRLyDgzOcuwDAjXOZDddCba7GnqHpn/v+cfHFecduvAYKaqvWdt6pAtBrdo
C1gHrLsp02wJkBbDPfDfyxs5qgI0ZAcyg2qUbgPQ2I16qbOQz+KHR9EyBXUq+O6A
NCx5ocFgW4p38IfJIPZsOtOPk8+ZrTb7bbyeg3zGDpxBQEQF6Wog0WpBPvUBeTYI
8ajbLNJzmTRYJtYwo3afMmmklcrqFPkL3GcVDM6PQlnl57siz6Ci8B46L4GNJr6D
WlGV2IrctVcrJbsRomO1VRckPlkHSwNqGlKV87MZK55+bGLNvXUDi7/dISFJSYTV
m2HHhQsWxvdkNb14tx6k5UODAg6eJsgvsuve3VG9FyE5rDexnVNc6ERfIb86FEJL
mfvyT6fkgThPa7OWAe69aqtSCNa67XwyhnBYELUzeRkLEjuC1dXIiZeSdWa7wd8x
Gy3Q2wt5YIn4KwCMu9X/9B9sLhCqApvuE39/vJXcp+Z/9Q90WU/RzTKXkpXUKy5A
7aJmsKlZVPoWbkd28JzVLvpPZcrpyhTJ714pnMp1aqdJeAK1o75Ko46cP1Gn/bkk
h1ZPC17tm1DrhOKFZnJW+Opj+0rMSrncN0TWgrejhxTOE04JXvbzkU/fiorqECgA
R+t8g1HexdNv/y5GJueS43jhWEJbk20LM1pxjUscVLPZwAT8iMgVtqZx0xoYqfwU
qDaShDBVp6vq6X0U39QoBbxKQHmSuG7gmabCs27bFTg+o0KnqqjUfuhiESdu0PXe
6ZrIXJjtnVE5KjBYUMdM1xrBuEqmp+7QkE9Agnzv1FxYknfIkASpGbxbrFieFXZJ
ee8wXvhV5oYsrTXDICo5qvRY9oGEb0qa9Dk2/KPFMYgakQXgDnYq9nPeWMFUl2PK
23WyFv/ccekOqYkmbCPmxQjMrzN1EpIusbT2OeN39hhMvmvkCCkMkTSBWkFOXyA2
m8jAdryuCC+vpYbnHKJHHZm1fuY0hKn3udfHk05dzaNnhjj5ET4/RvebZYGfNqXb
TIQkLoLqdvh9q1+0CQfIM4IUYipG7Tt+hQjK+QZhoKhY70LQvFlsuucwbJ8M43uQ
C/72bJ/i4F9siV24bbBUl6C76ozFlrzLd9O72CAcBpYTTFDZcbMihtN2sSmk7rzj
7sCWSl9TYr5GenI4H19K38xAys3WsKibIx+atjaF3pAR5cd00hRWY6I8I2JeYrME
0UdAbYtESlMWzM7A8i62lewEgUHjBZ3aboXuQ2BBISdFQ9yhUy8SJkpyU1aam+pA
OQ6zTdBTfFwXjNg+ObofqYAfVlOvvbrahpRM+0TN+9UNxON+mYwhFmELiAKlw1od
9W4FRk35m1RePbw6iXV1VY322S4pXnpM4wZQezHRBrNmsd2cRQMQxyR2PkyziFgY
O5FBHOXlx6ssu5/Ensb4SFF0zOBFgI9xBrDqopAvPtZrAqQVlO5Ilbi3VvFPFysD
p0e05NVK1d2YFSePaFvSa6a4jw2Ow8VHimgcCVpayWBZ0/HbLR3ve7f+yccr4fmN
6WyLJEIyoHV3io9on/UO6ADVib9U/Sg9XVT8UMFGk+DaofwylbQD+m/9R58ot3bn
aqKKo7mzRFvOf1065OznQjSGkM1jxo7uN/l7R1cDolsppLEa15mTqCtihAFm9r4L
T3Y13cLItXzgXAAJlQb2HScCu6pRAwFRe5PlF1PAg7Vy1kf3+vC0g+SsuWaaVylJ
PRMzp+iMo3elO2m90i228+a/bmsFDW2bEMmHgaKtAVqLXf9WyMg9sj0z7Yj0hgX8
bT2H6uy7mSFcY5LNTf88JODwheevL8JTuiW3tCRCJ9tbj+AgUJUtDUWCq91O53fZ
rZW2QqQOlsepR9FQcBWc1Cb4BH/rwhhTHKW9g0JFRwNWU2eO4kPmRKXaJfG1rEFK
Djzku0R9XGPhHSQcDQhsROSx4IY7f1iub4O2RSdgkuHPifvOtgchE2wbuIaJ2Uh9
JRsp5jz8iOSCk1VEsDBq0/8hwawjWH6mA6pPDm59TrtWg85h3hYleOBN6pWKRSsu
evw+AVe1r4HYKa9bDE2ZJqQYF6joZB4CjiD2QPoUYFl5sQpj1yCcq4w1oxGhFsjd
WFWBFEMNmFz5H4MFDDqRX0KnEOGDadZ1fubhkEdN6B0Z3cXXVpNWt8xSGlkUjpGm
wywimDdvtttNUpMu1bJRJL6qBYk7ORKDugI7znzfXLXERwXdZpHPtggu3ehKZgPV
8xeOvP45Uc1B7ntAS/WNpLXDy8NcoDkUvmfXkyKu25p7TaXPYV3YpmrxO1ize9DG
EgA/FC0BSfgHBr+eRIpwtVVvGLzU5IqWYOkIJTgNgRjfXFi0r7HJfc/9qnJbGzJm
PTwDRK7D6TjmX8r92BPbo3UQAKwU4duiENlCBLHwA4WLQhjGeBoz9rea1+rS3I1Y
2NllToJEiP0Ih2kyAJiaEz2kFcpqvxk7bzZGObZuPc0dS32fFBZV6aDltXNydW9B
DoZC74VF7xTDFqby647gWbdzlDeNouDVkzeWvV2r69gBnM+jdUhDOo04j1tlwlaz
wYgnw9Kc3S0J5LvWaFsSQzENmXgcWARRSTGvvONCHUrmYT+7i2D74zn16Z58mDh9
wjQjMZp5nDMlRkTxfdlss/jtag/sZjPsPgHDMtX7fh+rMTRBvhpGO0GfH24hKQsA
UTYRaXQOE6FzTRwVzFeNY2HniZX84xugvux/dh01stkdRwifXgR+X27JMZKcIsfJ
JsYbkTbxtWidm3WXxxy9cHE8+Ev9H1yLS91Dk06g76TssN5t94Zwdx+KfohmDJyu
NmBF7jFmoYoCmSBD1UTxkV6apPt9n8YkxEM+Dzol5tKEtDalvdwwmgm9Yxt9FmZd
AGD7HnQb+edV/dU+BN9+cXJXvFWnjBRZ4PR7oazDdIZ1BR1JbG9pej4MgfLcvw+/
a9tsqeZ3Loo3Nw/+PQco289VTYqN51auw1vzINujvfsm0XQjdVc0PoZOJumt8kQ1
b/UkSwyvu4ZevjFD3VIYQfHLGv4J0GE4NIPbvd1d7wwzbJp7eK5DT77J6TdLrYlS
+Sd91dgLFS0YuVHrQzleyPirKWG36ayNV/10NzlJ3yeXqMVQHesQUfeZqtbFLGUV
ntlqIkJYzHM8ptbMuPlTNzIpv5/7K6jxrILSBwxA1VjST8AA+Kp/s/7eh05RIt5r
qS1SwRbbAUo45j3Uy+UleRzqgNZ3QD06EaPoo92tEHWA89jIKFAFPkCqQVxz2p/G
ic5OxXNr66HSY3NBjyHJPWxbzdT5dA9cGStZc/cshgbpLrZhwpdG9N2eu4g0qdVC
9HlssBi62o9s74QNYNLqbBAmyG0z060fIlV9B9BXkdQyDt/Gd62fQuDKuZKb6mIW
elpBeIQYM+BPfsZIIUPbb8JQU13Du4rzE0vVMC/X6b0FAIoPA2w97OvrOF0/bY/2
GEUrLNofN0/pHJd2zWa+3P7Z0IjJqWuI+fzTy9gU10rvpD8DFOauTrrjE0bKyCFN
i3x9wNzebm4x7qrSVyjjC2TR8GK+qARdNyygUNZZNC2K58nBWkiTCUkWKi1FMZEN
D0KJqHngeVYLjdNanxwSKSnFOsLFoANzFFj0plcEkeoOxmC5Syji8I84zqbjZm4K
91Dkq5Z0WcpsBMm1eTICriB4okeA/NQNFMoNj+AUo8d+NFkBafIA2tJbzTySEg3q
OCz9Asc0+gUN/AzhqPuKe7uTx+5+LfrD6pAgsRisW1vkJElkk6TN8KfhZR7AIpTa
FIl0YFVvN3Zuy3kBCkgGrQKd03/T3N2zWUnDzDIvmIeRqZChHutf3q52d/5/WkJO
Hy6ODJgyWybjBpl0a6zEhVuZPP/Chi+QR3C4lp53dwWhcn6NFo9qrCrlt+VhD835
R6WzzJrabXOXlOxJIu+QPWN+ywFRtmQzKevxgEd78IYQJpoqhWgjjuijHa/aua7h
NDjvnrs5MBOpeiGjHdJsD6mJOzFpxTIBWxAL7COE/OJDaQeHxAyQYQHHa05u2p6a
YQ+cOzTaSgbO4of5xiYNQNjrwlGUSoEAmjO/sL13fkruo3oRm4lLb/En0fGOeB6t
neL2anqg0BO1NKFXz0XXwOx6RYIZZaIAd6D41NA8l3qgaTZ/S6RYVmYsJMq2adJD
mNTSCoQwcKGfj1NxMfZBos/LZXOcMzkllwkqBf3u6CSwgyEFyTXA68yGbJWNU58R
ZNo++nPeAccgJ6dfxjDcF2TTbYelFNh6qq8Nz/b65nqtR9cweaiMtETwgos2iysA
wSYK74fHgkspFR3D4cR7KyGlES+5Mfv3HZiN9lriKVTUkushB2RiMUtHkpG1I7/d
+VX3o1688Q3evu1Ir1AFBNxAWgs6O33E4/4ddR9JVMWOx4STsGcHw1Xp6hhef+mH
p+jks8Xob8A/ooKz+SyLmXJ40mx1BkyugdVIH9+a3ybirkom2i8rwctotIQG4LKZ
gDqwVwcjNCWwlATbc/kIR39GXBpBC01Y7pVsAutnmVlJAWV4pX39P0KyDhMDOXwH
IUdp2omNiO0VyN3CTIukjVoCXBChifVdLbtDkH+elg8ivS4/lz7S9N1EKppWPySb
LwMQZXdN39uC6mDGJZf8qqGrQ1zW0LlJtCXJGlWQ9XdTRYBe1OkGzk5Lv9a2CnnX
CQDlyku7VptUyNcpYQfdqfJ4pQXoHrarSAqCEz2DXIB1sAY1iHi4KawBoFqI5Bn3
7XKtl2ypESpQXlzd56dYsqvt6PH4Cp7kBJyH3hMGm588XD4JawAXUOzEKo0ngStE
36724TTwB0FOZQlaQrJZSJhBk5B0iHS7iXU+7YaXoxBs0tjBXSOcCBzzrLCwhmEC
6Qv2O99s1cvWsvIGpN5tsJQBU8/+qCC22KR/M2jTmK4kLiLBcqq7z+/KHjVecdZK
aZoU3JUeb+4jq3hVRsIqtFGIF47Ruy7EBnMvvkgIrLbjApE+MMs2myB1Ar7d7KcY
/px/+Wtie8TgLbn//datVcAyOTmz0x57GiqC3YxdeSNHzoAWrnEbdzKnpPgGBbj/
tP17EVJYp0QuUzn4uIIu2pakB8/Qf3zEgB+uk+DczYBu1bDH2slQcg4M5tZUiah+
bQVGYdHOerpCUttaeN0P+BC8GWf9hTcOjJ2741TJim/KApenVSD994bGPlgaXt0V
mJzvnJydFQLsdtEIHg5R/7Zq+uqjyLvnCgKenB5M0dhquqUHmjPugGEn1skpQN12
5OWLgHakYLZgczPKAUog7KyomOJ5q+5lIBNAhHtmDmrfEjkMOvstIezNBGYn5NsS
dL1Lj+uf8+QOPHda5bNLYoC8j4P68UQNseEI8DKeJatLJPenhpO1NBHQt1I69TDd
aceTt3NDyFcRti6DpuNpDUDfQoaGkwKnUQENdDXguCV7jzJLsVJTJk2XTFJvcf0+
00+eXnyCp7uPsmoE0A9EtWdvzCMGpULPuQNb32lWWSHL0HmxnJFhK3qBEbrhwsHZ
If7MRZPnn95sA/a2E7e6Iuf+gnGtyrFfOlSC7myMeBXMBHXujOBw8zhS3DCkwnk2
sUj3EPVl42E5K3fufLwthvziXRs74dr7wQ9Ok/Ma+jZ54r00Y4XRz7yBryHNiwh7
98rQ/wL9URzILut8uKUGEWy08sVS3yu0diI/tJh9JuUCQCUBZkfGQzrE5XlRrPGr
HQ1W7VBbn6hVqoCdQZMf4yuMg90MrL6qxJcUJNgEEgr35jXM/9HeVen9hXaKhWNp
S5QqNoLr189veBnWNnmPuRufTWYWjZqoIRWklXO7qzNc5IHaAQ2a926kFZi7Pl8R
zkt34JCJEFWpa7FpwvUz912Mmka4xmF2VJ8tp/YKAkcQg24UVZU6UxPPJpSY1HXc
g8Lanoir1/RGJUyPqH9jGfbYRdM9UZe4EL78CStSPDiBpI7eOxkc7U/493qVqns+
UwmyA/d4d+KeRCh6/bmxSX22b7KGT/qy5JLbENiC8SnUrRP8sPNfh+Fmqo13nJc7
0il83u/2R02laO0QgngFjDvcoCq9OH8NLWEpxqhwGjT92WTo5NERFIu0qV+SH6WC
rRAx+4Ui8774MZZCLQyGKBOz879APs/Tmpv1g8PodNg0b9qdJEaXeC3kFb5lOI+/
lCNX5Uxh3UxSCzIHvdrERu3pTmrZGycQbzJ1peo0z4biuBNGwMAZ8npQSfswgipa
q5Gb84VhrqmY9OF8r876LQNq0iIBGhfaPbtfO9FADx27nTYEyIOdW18Y/cOSwPZW
yQZl+m59n+G3HHpO8Uqpfv0cPZOUEDH33RXzwUbu7SieuSlQN0wuIQNOfzxQshXs
dlfSfAsl/ElS2ffCoMizDXOWMBimq9KO6R5H4UUQeb0Nq68roQfwPT3eznoDgc60
Fc6cL8rHQhmVTsLmtv5ox+v8/bBlUrlAeO2qclLajWHMGZXBqJtSdtz3ioUk7ZTA
QIZoP/D8lNoYap9HsasVHg3o4jBWShjXQ5Nr4esZBe58/hsMMiRHgxpa1vJ/NTuJ
mloGfkIMsd/KTsdcMo5pKN+fSgGLeQt/8qnraw0F0Tv3bZsXClGqMN8CUlowa/Md
va1jS9I6FLlMK3IpA79DB532CwZBnhgrHvE32d9Pe5I6gl1bA27U//T1xS/hPOLx
Miw8xql1Szir/KZRhIlZn0LjK1YtNutMTF1eHlgiCoidqlD04dgWi7SibpjbwYqe
iWbVpZTiPVjLj6UhKGODbKF2Qid/2d97U8IbeUW+/67MBi90/HEunCIBSy3GPbik
qpY8+aYqekpyrVdy35pPrwzXQiHU59ojHnwt2FrWpczqIIBa//pCaB7xWaTubxW/
ae3hMr4Q6nqg3eUJD18YG2/vFQovfm0lUOzBnbFl5DcJPIrbj01xLUCLP2QVDjUK
Fu8p3VfcedIXK8wDg6E9W98eggDFyxckc4oDMCyiRLczXmrEwZTor3LQ9HjqIIvG
Um9Dh7MRLNn3tslRqXmimonZG2iyZ7gq0obx1QSnaE70ZwTIzCROreSeOh54uWJu
WIOjW+tDl6gu43LZef+yCDs0Sgs4RYc/FOgbhAzAK4AudjhAW+eJ2yaaFeGEzZMi
HKTEuZz6zMaVKUAxVto2KbC3w1s9eq6LZK/IE57K2Q5Q1huGJ5CUFdmpnxvUclw+
0NmRX7LFQmKOKFcRCbHG0t8jGP/Tr2aZlV7w7fJMQVGqBO+rd4Nv19mZHxKy9wea
NrfWKIYmrbr0457Ro9tLGAdnH7YR2QuYqU6ZRCGqL4blVfs13dwMQLzo1lUimYqf
8deNpV2Q7dc74ChRxEzKuZRh+iN6KrSZh03a2ltTr5Lt5iBEBUucQDFcJ9TgN7Dq
QdjPGJOmjZmwyXmvrm9uwQHkhcOSP0jFHrDeuadqhH3wLgA3sRMbkTfNgzxQs0Ki
4s7Du62OgwgMDq5MZldlJPHd5ywvQm5czT9+5SyMdwZyMLHVElXg+AuVhXcq5hKZ
pYWb4Y9oh1SvDnUH5E2VDgd/bur4RBFlAj5+a2SZgdUpxyXDDsKqKMqQw22ImBaw
rWrbcpTa9iCrDP6i/RH/m9WOkXvwvTgXamd2oCN7kXzDZ5GNISFE23pvcc3lp140
vU6Kq/hve8/0b5B3mLG7aJQREh4sXPgJi9DUszOWsbothYxfNkipenGgovR15qjc
yOmnYky1vyH1mYqyI0lD2I7R5NKS/2T6evFNrP3oBBoH+G9n0x1dMIKEor++U7rT
MzySGweow1XmcP6Uu9JhVwf9tc51WX4vZQrOBN5RWIax9ncq9EtO13fJ6upD5sAU
aJIIqrO//YEimkZH3jYsKw4A9qyhd9U1clbRT6430qmaDLOV9XLywRDg6NrR/AaU
l2SfPRckC1llN1HI5rPrma2IzhvBwuW0FcRZsJEPJQfeTYRynzm4c2b9onvikQAJ
oUN94Hb5fucnTUokSThOCbkGhHTVamUGNspAXEpyydlGYwYw7ktGo4frm/Pkg9VI
dLUVnil36tUbqsZIv7Ci9mAr4NbOUVilWdwg+Dza67I8br3IvdR1GQVWNgdD8Dlz
ugIdXa0F7JtxiMTz7x/tQiX5YzfdpTV7V36YIMYSYyVpDupzfsoOTJMMw05g62Uu
N+yf2gk1sd8v3LRqUl+CRVRzghIvY1OyQDVclTK3i/na0xCjHoASs8Uk7cSuizJY
Ihr63sJzt1XJdU752Xzxqu+0FYSIr+3dZ+WCH+F4dxTwj466mpNcr5Dzk0ugN151
ZbUiPPTQ88DTWXJiKe2cYlSPuPq/or0PWH9s7hzy47cRFwkwaJnUVj+gaElTXP4H
gv/KkExG2HSf4j7QDpdUQiCGbpdwtLfSf8YCAVzJx0kP5y5flj8QJsUoOAhz7hq4
WClVPcSLcfkF/Bms+haAQS9fL/6eRsTs2/xsT40EpxPp/SWSnaBSUIV9kpPfOAsw
Xwz4w8YJDIe/ue7P8qmWMDeloKV5xEi01yrJmJNVt5AVBS9Cju/9Bgps2Cw9luya
fgZ+XbWsAaw2b1rFahvmGO8YFtHGVQdaM1OELiy5ce0RwLZJkcZamohVSRRDw755
VFZ+RJeIzolz4mY28rOXBxR5Vwr56YmEbPRSwaKoCf55pxnm3HCziGKFWgYXMyuF
fvoGlp9aTfweLSZDl6Ap9XfAC0nOr5d/3JGvHM1YMJeJGovmQvWBGKo6dADDXxdI
atFdbrFo6oafDufX5mYIUovrpUN5noklKt96uMO1UMqIXhDoj67+zQKSF3nVtOij
fPPlQgLd33xE7+v3siQE7qICtLb11l1ILPRXkhd1EHjZivLZ5oZ1kg/4agOAw8nd
5B7HIERVJlAOm2nnXssXN8P8TMT4n/g4tZk5MFtwAiT+jPVsz8x2II0th3lrCqLS
Aa9F/ZaluOYihKxUubbfTmc0Crqg3zv3OovEaLFhmn4YuRTxIHyvw2nzsNFO8z2T
ko4tsv9itjB5gHePo2cEPkXA5gqR5eZeeXMoRU42GUlskAjO3k9yoxjzfhY8RPU1
fcPXIzM5HjrRMwuT92BorRxh/8FLm1RblL8kBwLOl2wa8K5PTEvvdjRt0B0awzSJ
GcN1LJi8cGI8PZ50oyJKURgqhg96LUaiaRLg74zDRrsBpk7u5L+mc99bgtjNsY0c
2pqxbyttslayC9IXTXGDByouRCCB7lk6g533rwngHiE5yPav7KrNI8PK9i4mIwaD
EXkcuoUCy91yWwHeW8jrksfRo5HOcSoZ1BDFBQ/LN7iq37XdeXN+1LzMi2RW+u5d
rSwSKpMCZvOoPnfN1vBXUPtBrivMbAat0gPn9mwZFaMmwYYSqbaACKjgqJn+RCvC
Cbrf3fLCLaezHFTGFjK2g8XyeXbw0NDDQ0fSL0QpZGqXo32mfIZDR0e9EGo4GZcx
1hbqkR4TpKYH2ApSez8fyf1PUALblO+XMwtl1h/geer3jIwkZjarlyu2mK1U0gFG
1ebHJmovFZh2S88tevFZV3nJYM4n6OISEjL7/rkpqTz0FazuERQhoO/sWUXLu9vt
9OAEUhJR156gVAr3eobx1DdIT4q/pksfKHgdLHJSRT4XstiHusH49Y02t+8PrW4m
tgyEnc6ZBUBcVdWpZic4ybBjVyoWI2RLeEIsR/Dlm03hWBuY0or0U0dHuJD9zG62
KoHv9igVrXY5uUK7XBqSfhkGEohtNIPbEngO2bzoqdw9Q0p0Jjo6PEaF7l0b3GOU
t+8iTJfeG+fMwTlYJ0H+qCbQD/53ValZsIQIkuihwrRuSkGdQMVIKHHmsq+yHvyy
w5L8CXMVVfD/mHm/bxg30yqO6Tz4cY/z7IPuvB/7WT+b0Kic0CbpQ0MqiNqW2xdX
DNqDKEOy+giSaAtTZuVTBWYxdJzJduSzPTfY3xsAUCWFa1efvIBN2RCG9ntln/gQ
UyXfF2eRGD/nuMzEBlxOaAHPME7f8dZ/Y3mY+29+XNT3FGUccxxDC+HMjW9+k9XB
uxPIcoOq0DSQSTq6qcTRv33gRaxXmWvYvBXOOFp4vjG4DQrkfahvgslXt9yNpPPq
YtJdrmWw4Gzpyh8kcDFl+CBSCzYfy228eNVr/r9FS138xrXbOpQ/Mwk6R7tkRIH0
juYHNpAr9RgEfmARft0QRJmr/u45kFYR3iv7y+GKH0vDmwCSYrGICowQXg5BGtDJ
ZVvdgullxo12Xq8L7OrtsLLkM64HmHlBwvhoyULTdoJEEsslBlK2z4KnPbO8WWqm
RAhYL57Wye6HfxasdovDOZR1W0cFfiDc2DkUiSugp78XNG8DoZXUnEFzcEhESaZa
q/ijlwOxiQKC+Euhw6DOxc1xiy0bdQP+Kb8WUvI+FoSJGTeRAFHPxeqFjfn6ZsF+
5GkzWj7Ut/jj7uEmPdal2g9LqG8UFElEKWojyhFVdEvAYCQvGW6epo0tWO8sVcFT
uQn3M3/9FCGUr1Ow4beRlkc9ungxF/Qsmn0nDx9qHjsJ8T7lU+wISe8rS+/uZNdm
arzPpKacKtr+KEMyA97W2263p1GlDSfiWkE9AEmD9MHqz5SwobTGPsM5Dxv8LqlY
S4+iAOKrUurrEzyFyvW9bSkHh5WTfWc6j4PaZkMG+ejeC0QsoNMl4dTbN0lK33q7
ClJuXq16QJw4SCbmYJ7DecyFc8h6QBppdp8Px36K32ZlB6AedwsSP0AL1oISBCWT
sMXB8qwrzMxPsnUwv7vF7Mtx4ecPkS26uQH0dGpYAXzQ4AHbZ6fY+caTuCChsD3s
DhcPpyjLixYBRZ8k0bH3qXDpponj9AP3GBWxFv+bYCyk6Htkd20ZR+7OCD0Kcl3u
vP4zraqT/NNtwP0rWVPNsHJUrtzCzBOnwug2Pzpzp5rwZ9PTIx0/MXFneDQHae9y
bcCv7ij77VoPDxvQ7VrpqbmMaSPsM7RqXxHJMjWZz+wQw8KeSAnrjCaiZPPAmQ2Z
2Mu6lfZZTNz0lER2XrjEuCnkswlJcQIQGxrmWBG9EgQEIpo2WpxzED+BhrI8LHT4
1PAFq5PN3cYFfv9Nnpqdfp6VSeKWAMTKAjOIwugVE7gkmGn9gRrqjGN+OcHFqTNR
Z/QD6W1qLe+jMKqCrt4YWrfzGJnbKEYc0Rr4HrHy7u/7IW4kAgh3L9wUTlznkueh
27Rv/R24e9uxJ+KPgx9HOnuMW0rWy8Zs9IGJ0/dAShgtcytfjDcc2/g7wGDpBqE7
NlJM2ShMM0j4OnstcWvUoXeETyjmT4e3vO6XJWcb/FwKHkr1TYuBG6Fhkd7YBbFo
MUJYjhKL/ehkFVd4JwElBT5fpLkXTEKQ8VJmYWeK3M+SkiCYHWWLXsV6Ih+tuUAX
J/6GICfNONFb52+69ky24lBXp0PdqGNjDOxaY6U3cjxXyFcEfWg07t/oz6cyR2yM
bw1W3O1SBOrnWsNXI3pq2F49YuRb6q+yPkTSnMDjRvb1CrC+l5jDffQoycSjI9tC
MCO43jPzi8DC7JXaLd6zEdc/xanovvIv1DeLnqNxMbSnu7mflF2aLMVPW7JEsEEw
sbi35t9CalDkfYLRJOZza8R0TE/118A0SGjUZ7onm6Ehgyww0ur/rfE+VOFZJWmk
wLFIELh6E4V3sSBrG6g0H3fLPW1jQnTxbRRHnnyOx2uQhUwa5QNN36enbVCGJfkP
ZKjmHJ9lCfY0wDxvUslrIgB6XmmDhES6RwdhsfR7INUsXAuHyR6KGGY5c+hBMosd
yB1P4I66oLyZmNEeHMvtmEvhHbU9dlbgQD60CzuBl6d7OhDDIKBH2iFD+wAUX95W
xDkTa0S3CyzPou66Mc9/EKE7O58CNo14XGHkh4kAgin8K8oTSxIeRyTwL71TuBQr
tL+voiylRoAf24CO9ZVU5iz+wqkN+cWsTv3su0TdNbheFSyB/EHAV0vTe2MXL2ES
Y+Wj7G9Mfa/E/Ci9gSmyN0tuA3kckTDQZf8JF+Xb8yalS7h3Hv1Tso3cuaqxQynK
k3fCMCqoPIbfPK3D4OTG0Z/8XWp8FEOWHcm0L/jCPCrrnzy3BzLPg0Tmf6jGFU/N
Tm6kxyE89F+RgMWN4yEzmxu1fjxPxE5RxJl5tznmvNsQzAvEKD6fGwt74ttHbk3Q
CD4tvZiQ26VNgcH1PcO3TGvN3+VVKRV1lmEKbGg/6Bh1Ll/qus8ljGaMfpnUdyaj
yDgPfAjYgbjBU7RU1sGVTLRQ+tkLjhfaUY+Kgd+bD9cCNk2pXxa98cztsKG1r64X
wW60Vz7IYDPIlUUTpIl7ksTzei5IhNytrcli3ZJkP6OWsSNCjHpGoQrOdF4a/ckE
iAI294AlUmHwfuKUaz1JhTyzYZdzI83Fi87TMTkRgaE7f+X7efHWpTR9pd73KUKA
739RG1NVV0DmASO8fTcoLXsWe2nUPZGD0SyxxC+nFbM3xwLdJ2CzXnlbdi0nXbSn
ZsWl7w8w4j73FHETelA2yLrG3dJ9pdU3mNPbnGIJT+zVT7WN1tkVUtxAeN2V+rrP
Wfr8kYiiNPSBUVmTAoIt+JqB7ZUs31o8Onyy9M1F12oopQ+H85W1tZy6ZL9cxeqY
TAkePMfAMbPx5ULJl/oR807gK92gmEH6gfVI1fWG7pS20s50mdkIBRhdYf4rUq7F
KacW9MgrL97JjQfI4EAVOGIgoE7xv9x63opXz6v4pkn4i4c9h9w+GkqapjYuTxnp
yvhnPtB0mu2l06MRnw4KDULhYbSB/x/AiLl+wU+rjoDwWxm6tHtW6ubgTojeaQWF
iC/7dTdnJeikaDPPOt8vUWQgXT5LUEAMPa55oC0NPZAd+g4NPZVmZ/2NJOolizao
iZdpHAY8eAEWeJTtYWy6CsQ/Z3u4V0Dko6bu1qeLRXR7E/pBpkaloT1zF+xUS0s5
gB8MFrmuraS8qO/4YckDFGvuKdE01B8tLWcyK+FIdF2u81JA7Pd0YA6Leon7ze6m
PYLctRGbKe8p9q2zSjF+2q/ROmYzEgcSTYL5VMO4ZuMFLR4Vb/+C3gkOP4tTvlBW
v4HzE/PrSvlUCrtGqb8xQb+0T1/1SOaySfVmrsUwqM+TjJ5ezswYCAiaiT49mDHu
w+B/9r1S4YpzR3DL8eEyoYOUAV9dhMpH158Ylv3xWRyU0s6KMpNBvaC8MnskcR5N
rd4p+0qPXhSfdViO1U0r73i/cPwQj7MzZpC1a+Xo1EUxHe+8n38OpRlib5phgpRJ
oq2PHxqVzqHdvGHzJuveSwYBrDhJMGLxnwaSKB8P6tRsZ8oo3lyqbj2qQOE37WC5
tpG3mrUdSYsTg6QpTUfip3jSmz6cFsRZVnYbeT08JrYrwOFJweg20eobmcIjJ0uv
B80Ur23jOyFpvPTUwHb/YNQcAUpxMF0D4Uph75ZdJle470D2JakYuz0FmvfagVj9
TjFBoSeGkrsPUhuBPWM8W7I7GvMP5UFYgIeO3Q+sZYu/kfxTmQmb1C8R8z9sAi0J
4uCRoruCNpDY+Nb+2A+wg1a4SvrrdDCoxrCO546CiVSuxz46kuJVkcCow5NekHhO
ZIaRycDhwFmHaKpspaeX9DPQjuKnufRS1SilajZIJ8aii6IT+ZJLkicMRNppkY6E
TXWio6qDWvTbhtD7t/OohWJp4P0DQ52NCP9b/GSrsPmNeCwZm8ve4qkbvSdilhp3
/LTN+0f0cfUEeiDYLPC5Wxol3WeQG+gzLyNR4eHwCjIc3MI98eQtHVLb1W+lDoU2
VmrGFa7uzMcRzaCInnS/G/uKfUxywc2WGtSjTw1GcmxlfW/jcsD7v256tIGSKZtJ
DeZXqtvKm6udc3cfVgFF5SHVDwyJ33kYukUQwAtvTI5+jidMjlBdNsIryX60KDB4
iLdAOAurZ/2A2/HKYKBR2e1d3FF7jSM7ITCa2av2FrYFtlV/k29FDldNLBKJMm09
GKxYmd+shsUT3/Y+wmPyrfsVx4F7ERuSzKXaroRnVBSP1tnWbw+FDPbFjo9A10JS
FPVpaqlpQXUWAMWFmHdefFmKxL3heO+Lf80rNuxa/70nub1cbQCMWSd8b8vl1CUU
sYAoQL2Jg39t8VvoUb8Z+lQdGhFhNz4rhi5f52zFYAjFM/FRuWAn01Fe8dwpBTKu
WKxMlBCqDgwnOMxal9PQd1L4KKLbDSs9Z/7hQ6995VKs/NB3XcMpFCnm643uUaj8
AuKooG4gFviDYnBIZcwA+OVmGLLHc92ih9vfOCTgcNJf2DEctoXBW8bynSrgLqeC
7dMZ5r65DriT6yqI4+EnlepUb/DZJC8Jtz36PYxWEI7oFlvjReq8etiMo97kddsE
5DGIJW1Kn6/w7UIbUe6fzyMOXuCi4ZV3wriCOMm+TWf2/n9STowBrq6f0m+lNcY4
Lklnhp/Ui1g/QakGgkJkS7xOZsPLXWqOej4lGcEyeWUkOyoyKebYFdW8worpMxx8
3y4kEwvjw8/hZpHoAIhs2dKSH1tZM7YBu4ExkgZn2S49i+9Hg5SGZ3Cv4vD7Jfms
FvsF6EEdX9bS9w0BlgUgn0lYz2yvpOqxB1Mi+MCTZuhlQJ5LJyFk8XzwjSrgFZBG
x2EFmXo/GwCNRWPKxrq5swbV+wyX0I0QLoxsQxbIdlQ/3MCUZ6nBFQos2K75ww6u
EgftSaRhMYc7z9HfOyNtn73m1D6BAYZObulVsrA9LIWFbjfm+Fjs47vAn8AuKs/P
xkdGfNc5zj1pfMN1gKMRcpd/Or1p98AdTey8SwbtuOBc8jrvAqTt2PezMrUkb/6C
qWp2EPSk8RDsY1jpZ9ZERdajP2foqIwkwFJj64ajQ86rBbZASx1nV/swXtYd8Hwm
z03iM4cI3KlDca0yV+gyJzi6qcDWF56BOVLq2I0sbOk4Sfnz5wbkLcQwI9HGhv8r
zthvcOvJXuo57b5vmElYZTDucWmxxu8iNlN1vtY/JPkMxA4LSuRxBRDUbRHPyVmh
lC7G0U7SMQYSzD/tpz86YfK7DqSXFsVZSqripTB9b/lWWrRSpoVbjyoew8GNZOs+
6p21tsNYi9ju/nh/vrnv8p+9Moi4azElfganM4u878nJxesqZS6MD/nAyBqqko3B
lHNxdCWOp1J/4nTMhYIl14wRIF0zUDDT0TIQIi0WPwwjLpCOx5+vse/bmuBEE835
XO9pE+3DMvdi0F9KbOM8r7TzqLu8DECtcH+Uhqu5pzIyeh9yAkmclCvXyMiaQtMU
up0WJGTpySyaESA4u4Am+qaYpGkUZs2jgVfOGGnhJxgw2En7Jfqv8E7EKwBV+6kR
VP2QDsBnnsC32Ce7RHwM+FsDb793HA2JSfSEZQUsAW2v05mdO7D4rXdTlj5l1Fyg
kS1jA/vBkTHGnod++V1SQbkXAwD7UK9ebKBGayTHAZaSSYeX2kSDabedFCvN85AI
/6LxdBsK3TTLTJBWMKiJiwFlHpIOo2Bh7W7fqjI643umNWnxs8DICzQdw9iYAdR8
t4qtfFa7fqUnIqMR16h9Rb5TcnDthA59z92swvVLjnoznBEom1OE9zRXMwsnUhDZ
5aduWZupjLrNARWZmKULPobjfN6OsHL1NDzr9x4H2U5r866kojkd/TPYekAmTGLn
bKKyBRpHWqH96Xtkf5szE21o6F33aMaiRKw9sR1GxJW/VZT+hunhkxIk7zrYQdPg
SI0hfAubPGpEQAyAlUfy7lc6pE9XtIhUrcNsv3uQFXZp6r9N3sXb+9/Arcas06tp
ofTTd6MhyuQ/x12etGuizHot+U+ucVYc9Y+GjcsLdEQSGzjGCF8VxO/zOBeuBC8N
TXs7+3C/BZJtUHO1Wr6Xmrwnn3AWjvADE7fs0LAIS7+NN21DcJGhzvdz56YPu03g
vWX8LpQNtDUIcHRghlVq05ObpShDED+uznOCCh2i+GPiB3DCY26k4gjaQL/RI1ip
qZIiJ8pDryFqXicheI6WXhscThcaTX1FSPzPWgY3Pj8qYo3OeQF2qY3J0Gjf6p+v
1giYnaM/eH4Eny02+F2sTB4QM1//xoQYDIkg5goETeN4RGDCY0ag42DBLiVayBNV
h+RxEqblIfg9Kjr3yy6JLae7GtaleCyHioVsViq4UlSg5l51+TRUxRObF0H+dzM4
zJoV8Gg7AVzcz3vP+SDEDsiFKizHQkgZ6KZBlhMZZ3O8FAl7jofKfbOrSPgQsfUa
IOJrRdGi0Q1WWk2VyoKycmziopoR0bZ2OL33N96BMO/uyVKrlyOivfwLMTn+w0NT
KrHPi9YfyonK/uqDqpSwdpyTm8cbgXpC695+QgTNVg8QuOfHlLRdWz+98MbZ23r0
9Tqb2sqmzCuoaNt3WKQL/1xR9LQulL7CNuSsUXQkaNYpviw6c8/tAfMymQcqWLjl
9fATFOCgMxdykxZEZrvcDrcTBx7lQ5IJmVVjprji1Mo81ZtWRn1HKMOz65kzw4o6
VLqPjVdi2eoqZgyFwwTmp0AWzU8gpCHaYaGsiGGg7dio0tuTDNyh68hqL+fvzBq0
a7BB1ZiKAOwv5TJJCamFYbCwiav/sIY2kAOto5yqOsFQxxfypNwlRfbfbKFugpRB
/QEm7dTsecf39INFBKbDvCrjvf90rictXxuzbVb0rJJnhF/TGWYM4T7C7c3YiavB
SKcCB7xBcVMCV6fCg07NedVPUI3JDLwbes0CRDR+KMcxd4DAzoGJQHpqOyVKuoyq
BpHlobC77MzxLZDdtijbD67h/sGrKSXQkj4kwzeks8n1Pjv2+3dKEsXnLEWdnu/8
n5fvKzEk64DtY/QyFXBBUbIKMF43ehKeupPPMf9Y66kQkZ6BhRg+YV4EZKRFYyrZ
vEirPWl+STzm8upwcoBf0jKXM3FQ+7CbOoRI5N2rgK63p5PfT3+YiuL1GyeCtYbi
2Aw9Z7b8cU6OPbCD/cpui1IxYzoKIB5+KXlpeb4n5ng4mjikhc+Ws41zvqUXfeQp
VHyYArdDfGcAjKTw/vw2IOyxTDjwXwuuq+0JYjcrX5n+XzY7q196Fs7xaSrvrmjX
w0WNEZZd11FQlD6Y4ZYzMajn8kRU3RxBSm2z28Q2a5eU67MhfF7TWa5vKYP+5P1x
po0kjp9nnsCtFal8Q8MFJxVhG5ocEj/tww5mlMB8pdb05DfaiB43qfHdbr83iwPY
AUYmVd/RU7aRuJFDue6jo0pEPOzyHNmsfwURCCohev42j/SAMEIVPnr/Dv3eJtMh
HjKORgw1zsRiDbYeFRBG60dodS+GGhWePFWul9jxezBRJVzrrmpDgI+ifRM3eKyE
ZP9CtOHSPU/nyfYI/cZGFVd8S2lgG3vOHk4hM/LNniMP870tv69NhBj0ibnAScxd
IWjOFKrLBQHD3iBa7BSe42q+OzpH8czsWU8v+gVBFNAcoHdYBXzefRe33hJL/XCx
2wFjlvDTUYs71/B4mWNNbk5+b8o8JA2j8bPp/SaLdI3O/Z2BXGgecAg/h/btpvPD
V6TXo7DNcPsEY9e9zFNX0S7+a8w7PkqpKKSt9VxtzJt9hZzCeujxRe4Gu8aij5Q/
Y3D9sPkaFS5Ig4i5rZ4IODgvNeuefCEdBLvglVd1KVJAB3keHmvsxYgpLZxMuWxe
TsmaUiNgT2DZffQ/7Vii0ru5OcLalqQle7kPPt2NZ4w7NaA6zegj8EOnc610gNkM
oW33urJgMlDLg3hkpK72SfDdzbsNcTlLVFg234V/uPU9HiKnV2rGgc19KyrWQVsl
2QNyGKsOSEydHrCqO+d6nb/syqVvhXb8SuRXXOcUGqaPBY9pKfOwk4WVuuxfE7dp
eiHxXNzAH9Yhv0vVZ7cuevNp045+DXRd+A1Ef35w5abqF6S9nvFQYdgmqo3PAim8
3BnFaVl+mINbzgi7mB1Fo5qFqO+D4x2StDzlxJGK4k6UBohN9qQ4YDSrFWvW6hFL
N3GhTxv0pAo5xc/CyaUKRCS4SFOGB18amJGTiZUGXBNgbloueSYWmSN/OTYVmj2B
zBbikMjJm2PE7LJ9UwvECazmFvIkn7BAZdb5cGFXH+CgW4zrv0LykujNeAqOypX+
4xS6tyWmdawYZK3Ke7mQsRTsShaXXjSVH9i7T92Y3n5cWyNZG5/mwf3MnQggY3o6
4G5erHICTMrt8Pv+MFttnG1v6hUpFN4eWEA7Av3VJ9/x92pKiL2EbPLgOx5fImCE
EmQ/Pv8RQT9ql7jaSi0YHz0EDohykQUOwDo+VCnMidaNaiivEpAoEOiEXcK0EE4j
aPP3/AI+ydn0dXNx4W2t9kzoLtozQkPiNM+mLwkL2KY2Ky7nbDv1QzOIrsS9VOZx
D1VDQ7qffPY6ZDASq9nR+1gykkoeDk23dvuvIgG2J8PYdshjfxhNLN2+aF8xyQGt
ZoC5wffHPukU03srpwmYq3GE6Axp9QlFEGmEh/6DxHp77/dqbteIFWglInSvGJyX
O8NVMGv4CWqC/xoIq1tDC1CyuzXPEvpDWb5+Lr2uKx38hbS5tkgwcGNPHfuIlh5B
RrUTssq0v/167ReJNi9JECHd2XMId5ouhv4gU1f6dt3+5WLgPnWpHJ/39x/4vWCx
5yze07aunYw+3WdMOXCA/N/8Y0V6vEaKJNADMGOM+i3BB+X3PYcujFGwY+a+cCmW
kRcPi6UMCcjI0qqlUaJZpcjXhL0jorFb3KDmmaOAxgsLn8FdLTqQhPj92SiRH1ll
ETmGgz3fioRXCVBcUhfpFIQQpinOLJ+LnwjFrpBAd8Ljikxo9SHZtweGDCfmVffd
NpAVy5p6wxxb84C7TRAsijlaSMjbyhUE2AulkVxAFu+aui5udf1SyWRKdHBEKix0
VArrWPEUhYkwqnUWoRUFUfzsiejqJ6O6E8oTCQR6baTlP4HUXsLz5BTWRsduZcHW
RnpJhHoMZjRXX6jQ1rLReZ0MJfez6nTLAcEPu+tYcRA3ykd9zsqVLnx33X5r8qqz
+p2c09rAXQHE/qZCKe67EKPBrmZ2IsKh+hVCSRUTU/djJgfUWe+nS9kUnfMeelYx
ujPLQNrIM9gjdwBIbkHnlbe+cuNxWvwSk7rxFDerwee/X8EK2eq8Kiw9ZaZMpYb9
61vif2eyzGTswrbtyqDFp67ZQuwoE8Vsv4C+SER31NizSYsIV5VQ0eG2d9kEyMtI
aJauPDCEbXZ+dLm7d0sFtwGKDlwarDjyPx3ERtWyXgKJ4ihRTnEH66KAEaxt6umM
gi66msm3qrbCRJmFvJagnKrMejDKCIwN3TfSvzn6NNKREcmd2y6qJWh5bkVAMgmL
dcMuPqVLftD5dJaXWf+Nwt/ztOUPEtQW4EdgxHBbqid31rSzIUsDmLL47oEm8Dpv
rnopjeTZcWdSU7YokY+tkEhMEJN9SQxxUbzd2v+RWVPQtYk6dSKGLMrSAPPYfUgU
voTworkIEyKotbOohNzrtSI6DKJFl3OZKcXkoNrexRVHxYbJvo+DKGLXaC2fVf0B
554Nd1/u1wkVzYuiVHcdBB2So8HUSxgVt6Mt7j/AyUDZjvi6AOJy5ZHEIl+sKntk
3szY5Ql69PXy8x614n7CmrTGwwm4MdvIrLG4VvEelSxsK51QtThJlm9KyE+QEBL4
VM0sjr6h3tXfIHlV7HaJGYxYESPPIrXFock6HnM9cTHHl9Gc7US/3CKq1baf0hKu
MmGKUIzTHTkJ3tKErQyiuaRtQmbHNHSW6t0+Jb+EWyDj5n8NlOaOJZAkMStr5f/w
fLdLQNVx4qZN/MQJpiXu7TgF2oI6f7gd7Q6Ne9LrfNvAl9t4nSpGI1pZYn3OJ+Tf
CaoVSuNssY/n14Er3+9l1VCkdJ0QLzZ0oevFvZaw2dzslg1uWeCbAoeptS1cCJzl
cvC7ohceW6iQRy8X93gpNjR1ValcbsR2FWgVmHcJWHPBZC9U8HeTaEV+dfys2vkF
uIrutGwiaja46oIx8+WRxisVs2eJGGGX9/C0Ns0TUKhd9cUCGH8418NudSR9HJGy
kbXncDBxL73zWgIm7ihEIlR5xaRTpfMnjRU8w4FYwCZ36LlMt+8+Kt+yGippEg8z
SEz/NreaTEG5o4IoJCzWlcK2xsDVHItrvzrUQhMhYnftLINzkTU3+ePMm/AdTzs5
1BP4l/E4hMvNjr79YjA7Jl9aFOcMr/w+J8zKwIF4B46cXnRK9QRzExBPDRwuPiT5
sZLKTGOzJbYoQ1H08vZhtQkVGFy7LJwEVltEfFouDJ317Mq0Xf0SLqhyrVMaaQOH
QNMhbKTmUJ09D9cNlIHi4NJ6JyGDPGzPeH+yLE9OtVm8KdlcziF3RgpttVFl7aSU
BdE6KbNYBdFcFX1z3mEbcaU66TSemwkdUoUAqmf/JpdQwcWBqsvtBVXHwYk9p13w
hik5o9RtjZa8DD/DhYe5MLSgVCOhxOno00+ywlRf8+1xjgliipraomT44jN4/Nmn
8oiOHseTVJ3N+wLepzjX2qUM4a4dBBf6nXBZuwtSqNg1+R/RP2qYx9Ak4ICxoG2u
J6FQI73bonQ1u8tUPFHJTxw6IxC3paFpg53wJmf7Kvxt/aFWmaKFCx3YI9FIkXL2
8KpT0D2g2JumSF11lm8zxSreudqlL8B4RyiKbk2xlI6qGQCTK/AVOkF5K6/Z0YpI
apR2R/Yyb1u/E6w7mgt0QdWiPVCi/9TbVPxCrQYCc+pNJ+bfv56sP/0ffyAqT33E
NQcFDmr5HzpMGU82eEwP8XhBPsyiA51RJINtaEpq7fS5Jg6bYDYb8rtJV1fW4RhM
0NM+U4aO5N1+GB9bNp/p5yjfddUfZvCFwdX5QuMF2BLs3Z2UDoZwRl20kJbNy/1A
Ke6chm2OMIQ4byeF+bP7MDWuJGUh8YAru7z8Z2g9uNOKZ/znubwWw5lRJBGNjcxw
/BIkPufRkt+cBfkKiSezOINgJEMUEhE0BFJfuOK259VFjppOSrVlc4m+poBbaSUt
c4vDWM8r175rbPrJ84nh9eUVHEXfHRb7f9OYsQ4b9q8ckBkarDdgMz5vRBtZ3CYI
UB9dmha2hfAaoDBFe0LtAVo9fzrWbzioav//XK3xN15ZjfS8lN1dbvouYVGL6nUN
TbyM2rHHgakNFW+yPX/p/rtrt5F7aCca4z5z+LoivdIpijvGO4LUI54xCZWaKEZX
NbPxYILOz59pctEgn5A2kTqnBometkpVdrX2US0+mV21HL2MNSVl8CP5eA9S3zHS
CeH7geMBMM80guvGmujunTGz+C5Ps9dCGAkX0d0wV1eQv3GM1G4C4mnBdBMCMGcY
UfkuhrRWALV9S3Ttt6ubtEujYE4u8X9mknKiVDU3km+zCf0lK2wUelKMwqjl5wKt
9/zMOYJBTpWHbZ1Yv2YrMIMavAy4RhMklVB6OkEtz5YZVRq41Sdl5f6KEzSnS9X+
xvbw2WmRkdQMFsJsdp/WVeJOHsJq6vAef6mxfnFc3tD9TpLXwwgOPNpNqagwWMb/
d/MrPXTqX+gwDYs0V/aAu25nWBYXUWUIYjmIjDpu7RpV0BT/kS4hV1eDFn1JvCFE
1U0n3pMl+a5LWXlNXXx4Ne8dYiovOYdOtuB5iNhQUfAVUJGnkwDCwbGmcatoIL7Z
3v5sFkBgdeHIMLmDrtMkoGYrK5Bd6scQMr3+U/NhQo+P+dV8MReHboBNAEZ7DPYl
LmV/chAPDcZOcsz7HeZ9xJsrou3WHeQlg6DWTGLLH0uWoacNnjIYkKGam2jHpfGQ
6xVjUtcp1HsYKiMSlQ+SIvLqAyRXVXX1jClZhBO7p14zyM8qPntaQjr4v7riSHpp
LJVP1S94FvQZ7OQjZ4hUOF03z9aWr2/1Pfuf1VEYIz7miSYm5vPISSOKCb/RMb2M
7QTGxNBccZGRVnC7EXe/DOJ/0o5TaQYWon8U+pXSfQH9bMCfQ+noG7S0l/7NsZfq
hQJYzJyZhKZl0uY8oj33Qi6WwN96KJHg6yD11AEd9YeLrySK80Xzyv+N5NWcwyOi
v7XwpeP7JYDyCGo4BEMmrhAYUQEZY6aYC9gDdgUlRA/4gpDCSuLi/65kKPu2xKa+
v1z/Srwffz7cSiy1LGTAWIBMMyXxaxWL9wkiIwgTCLCAkWoI+Hp+zJVamXo9I3y0
+NGASUEa8Wsce7BBWBdFvYeP/fQZN9gBQiGEVI39ebHqDhTVB53gV5AbHFNs36JY
IzdTPopPAcff1/4I1IMFn+JPATCwiypazsWm/4HvMCd8TUvxAxaNe5LAE4PY5J8p
H1v04uxcz5hNqBgrL4PMQOaUsy7F2S4cYQ9H1Ke7KsyCJSaL3n6iGVp/E8pnoXuf
hVTYTb+89MOZDhWoRHMEaSELdfc/vnrioDHEsNIJ9DfsP4WbSJwUJnLHP9ZeN6E5
5qt/LhM4VlFIGVMIr2DvJScSEkI6zIpmSg03wC+6YdNV4wM6a6QydOyJCLdsIIpY
vEQL7FiSLKxCdv9sl21mb492UhBm8CNCn9Nq2/fuh0CaSRQvNzaJxbs4J4ASOGf9
B+uOG5zDmXfmIu4x4LJPOqTqzQ92RsY6UYIFyzMlS8bt+mjmzNbQ1TlUK6GnCcl7
gAcPxBQvJz/HSsYG2KueKMzo0fpbpFBqtz2SUPoCAkaObtAEl1EWR/2n8e8lkGQq
jS2C5MxGsG5c0fDFVbp7kXlnDSldHi1BjFaJrP9w9N5W1V9vZ3sOhbqPg9sRqwhM
VbLHicJmIWJXHx5dDJOn7NItupcC7QAlXNlLPvKpjwSfZVaskOMawlFZ/sEi3pOI
jI+oYafFBPuh+V5eV1snfydhG3+uDdArsENNQt1QXMsdYFpF820+f95nzxW8//E8
6a2k9nJUSaH+C2J8734IudxPDYvQVEz8dm7D6Nu6e7nKlv/2IdluPlILE0wjAD1x
Ot+y9Kg22UPguZ3pdKwk8bjEZUZm1m9HcPDBht4YGJiqvMAQ/v2ceiSm/XfqQC7P
xb6x2wPu/7z1Ysy5n+ndAdyFdsRkx78S2C0OYF5Msabuz5euiy35GgomV8D9n+ZP
wGf1+1hSXQLNXyRHlCzv2IDU0P7AZG3Wm9Ox+5v2T5CeoiX39BXRYRAhX88me16h
dVRcbjyRv6PISEc+HeQffAQwiTVwPsmi9uK+lcl1a0EPFrEMSHdLN0RoLpnKY+l8
xoJ8YWIRzQcIi24J9eUZp3vbztUEYZwjkE7m+mV3dXr98PI14oQ/vGBmQ5Jn6PYt
GiwBGTbb0xwLYHR4dI/RBkoCaJIoK9xpsJo0jl0skZDBbZ5xyGPbOU9S8FTWE2Bb
47roIokM1g/8nwEknrg1MO9QgI3WazdIlrOxXKSLJOOtojQBJyFcKwFaylq3KOGP
5fYe4GYoOUdWEE//6RL2OYYQTFY4+SM/Qd8dMpF9hUjZyC15EEQ0XFsaMwrG+O3P
woBBuQD4MX+r546L2PeYcP5OxgvrLeYN3sCuZ5xz8EDVRsc+x3uDfoRtplRC7YmM
eTLfv3NJO7c4464za/hYm3ideMLnIDyVwneQRrwkM3BCrfyjkXX5ObNDgL1lTcEP
XuRRY43Ac1jY0IDeUTmTYjctPuaWuEut6tZo9YaeOY4KbxstcfQRsph8jKLdJr7n
lAFFgOvgtnktfKxPtAr6zDS4LTWJpT1gCFwBEiGyf+1ehLsT8Hb9uYW3rm4MWZia
heNOFDP/YP/nTDEixLpz35l4j0nNqYjqzKxEGnA8gEW8qY7nKRj9RSVrcZb8WGgk
xH2DVnMXIu2nV956as8ucEGvUE+pngIHKNvhtb14gJ4gdvfhrh+b1GaJtD98fm6Z
70ZQprW5z6bZdmvPY8M23kycjTGi/TB5Myfh5CKmNzoqn+cl/NJorF2XW/dh++yb
FuBL9W/THSsyBvj3BjuSITD+lKsOVX8fal4jIiYdq0dBbOjMLiJOQdwTQa826xlk
nZ/Ewg4+bcmHRlYoV4grerMDAISRK2g2xx30HILUVmxZBKFaBifGPJilVz7qEMri
E6mUvQD1L3I3DD9Kngz7GmLromM4JltxNfB8dkpz0teqDcb9N9mvEYOy7+XZy3Sx
hyP1CqR/t9qjnD0TkjivVdKSd1AcKsie0wUYkvVJeXZh3Dq6b5JVmS9BkyRLmgDT
IlFzSKlnUnDaJmx40jOIR/WIXp35l4Iykds8HN0YsEygbMHJfms+89ziemkjpHtd
O/2ELBNZpn+NAAbTpbXauHGeLPteURcTfYXbCl3cAGXry9p8O3SnASmOLwF2Ef1Y
ClsS6VGKrNl9/kH7/6k+t+hm086fQTwa9yk4C3kkT+TBEQcdcSxo5akC4kgQCzxj
2N3wu8UI67kNiONzf4RRYcbOARuXsTbH+b3GnlC36w51TnpTx/NJUM0pYErkzA3n
0WNklcjg2JWeIPFA0qJqlFR5+pfL99yyQCYZr1e6Gfn2xBbre0X3rzXKk18kr7OY
30lTERnsDJDI9EQtoSkt3RhVI5v9FXIkLnoxTpY3VbErDH1RUy3im/h/qT46Elhp
XXf4IOqi2dCXeo4arWJKzwe7//VgQ4DZxhQuC6WJA5lKz6D5glsNFZ16q5gwm6xD
0tor4ymcNPFIFOOHfUT1E5GEbB0lFKZ0QyaSENh/UtFD8VbyKzmdpZaj5SKYSh3p
8DOTxpXXIkQQpaktHGFoXOod8HRrmJl7dOQXkw7AYq9Udvs7HDIYh9isUhjZU+G7
UgUVaYD+VVGV/zy8iTPGAKNNt3bmS0U9P4qT3dGO5EAlQ6RE+CKXHPTaE14vushe
hsvpJT2ZPARAXfECFkOhSL7C9k1c4wIFRs0ybIewDGiVUv6d+46YhvTkDMBBKBS8
adDiEa1YDgKtBoOZzJbyb/XCc8yXJWDYUOX4PU/haAR2pG8lpykPrmWO70d1m9yV
mG5MQBLT8Htqod4MNLeVC3jQ8Vzt5ltBTdHsN6WA94ZmH2jN/B/aNpvLhKTvgYhH
KRfC/w8OHCV9cj3j5bQrrzTwJGj1uCZwZU+gz9vHjvaO2SryPTJEjazMOhx/FJq0
b/u9bUAr13eYSmJt+k0ffXfWS10Yyc00fYnzcO4PJarvN1XUkRVPHntOiDovag4N
bLogNebwDDqZcbG5yEewr0XuhDDqZ51e5RPG9fMw7JnVUWD/rNuqUDdOvyFJFYxn
+O70XCxMzCZZ6biginFeivN+gm/CxOBehDN1KSbSrbu7+OcJaU2KQezfl4DZMqbk
6hZKI3aPAeeEeFTwE2NIvy8lEXBEV1PAkENwdRoDX3hmk8Eg9exiRwUg2wfPunaT
MvOeywk+nrlb+Kh24L1uT8NbncCm228qYqHsn/NxkyyQqKqLOvBrVx/C70I5ed0z
982IsWMyt0bILZazd+SkL2ebERubzxBBoQbxSZxk5CA/NRT2lRkGhfh8hN1bpnul
802HVscXbJYAYrvM0dtU/jYYBDRCCsMLkEKmNScgzvXe8VfPPVVWK6FRVJ56KsIU
S8Yn6lnJaSGSUvWbTddEjOykgCCreQ6QEzDOtw6NzTgxS7yzH2L1xO4aTfCwoAGq
lKI4JO/8RVYDzBcKELnSNdQgzLXzJyanMruI0npLmE2QQ7g1+VJWcWmWS6dU9kDW
OmRPDCWcwrKABBo6WZdi+nW2l4d86gq9tKlQRuRPZ6txQw4h1EYrBXY/9DFDG6uY
15mIIyTgO/QpICD469pF1R/GKu0vSNwbUJ/NpXeie0enOVIQs0sZdRqGEe9zkkmr
OnQREpAHQpyF+rwAP9doLFVCroxn1H9mMstHNysGGNSLAQioB5nvoqcbmtL35EUA
PmEnZtusCz9UsY9xQkqz8AwieZT++rzeSseFwBvtCo8OiFDAhV1ZokJz/qXeNc+Y
ukbziBOE9rcOPttMIlM7oeY/88h2xgFo7YlQnMuB8tF98s2NUly5CJ4qrtVIaIM9
SVyMrNvqFaocSc9BMWV6fFlhnwZdjXApNjE9eQe0RzlauaUIuKYPZdHohCkyW72I
jMbtDIrASxQjgxQerPSUZBECVzCjhKxmJuS1Yb5JYOiXgSEkOWG2DErTcOdmWh1S
/cC6ZRGv/YxZKwcrhp+Mu1Gv+fqzEZNsxAbempP6u6EcATzykrWNfHXAdqvSJ6YA
TjGpW5XyC/G6acI91QNhLgvQg5X+vD6AwG5F0fUHrOL0VtqPcHN3JFRdBZhyq3pL
az8lEGBlqKPlqVgpg6gVL7b4BrSmUMFBx/m0UtRbQvGudbCeKRBUKShiA02eAxqm
aSCpneNZIxMPCn5wTBWiffe+x58y8YEWzQaxK8LDlofMciiUm3Gi5t7iQHsp2Ahg
FoSTj2sEP48VUcrHtTG2o9P1dETcptna34if/tqIZkZAhsj1qTZynQEqJVQTM3Oz
W7AheNS4LfT6m5fHPKfxaWiCsRkptay0Pbixxqh3hdSPiM78RnFfhYs9wyg+37QG
a9zaQepxVJjNY16dNkjHoQ3ZsSJ7HYItNfIPlnvxyAJIDluQOkU72JIPtooMilYk
GlqqSDxgjOTMt960tU+AhtcxZnN7s3yEcUpWya/tT36fkTbNjOHnBxEmpuG49sX2
cqCHcT/9CcvGCiXSErprQs1sjEDjFYa+UOHHLJreZsR76XNBM2YjOUp7enaoamCA
S1fda+h/Z9XqAQOAK89zjd8B35Nqal+TkmKSrKRysqJaba/4+z9/uJ8HDPTNgxcX
ZbX9R28MN15uFoQ5mXWVaHiUbNJNCcI2pDipTzSP8x7JFHlAvMwr9geYcw9lhLnl
VArFSyuw1qnUIdYq9As8Lh/qpG+JCwkkuSQJu8Moddy64y5wMWwXOlNAy58fmeo6
Y/evK3zYjmCAX4LEdevaTkbhzKw8FzCl1pgjpiWNt+FDioQ9g8+OsB7dDdPMeIoK
pq6Dx3+AGmtqciYBxQewPnVHVjquwIU5RAeZa9enfJXB7QCwrgbl0iRu/N0cn9B3
+8bvhchmVjAllAqu81etzelOtQ6wL8pVUBzdJzTifpzpF2VO7645+2FNu+39W4z8
xy1TtDqmMFCCmcCMBrD9bqF7sKM0HqBhY8ESjZFTuJrvjVBkka+zHx0we0h42c5C
tFGq1K7JXhq/PiqWx3s6kz6t9xmuMFmEC9QdHKHoBY+NxgQNNTjZV4n5EkquqnqM
dj9k5wvgkDjWb5KaWzmzNjcUcb3ZF9cKAzeGIYEkXc4/RrLoj4WPbKuvjVaK0Vut
VaR5bivxk/Ai8nEXmnZq0SZATvbTU3wk74SLJ8pdQviY/OwinS50gUM0BJ1VmUZk
h7M0voj01qlXeRhO54tMiiH+DJoNVeQ4wrNAuqboITeXg8aH/mqRxuksU1LmvbMo
YNs5akP6yR3w40899izTeyC69nXhb4Gc3PFplsYkyRfXw2dDIc+bKHRulRQjk+Gq
DhQbqD1pZ2utRJjEVXryVtMHLuo1ApgZVadhyHJHHH6D1YhQSfLMdVhyzpu2uPEM
DxCuimFaXeUtvapqXCFu1eezpo4XnsPWMFHJ6Iy0Km7yH8K+D8YbTe3Us7VPrcuC
hNbJJUZlrhltjZB9a0nOG3tG2YgPQQvB20IDeGsxdfnHmdKCrny212zqjdB9aJ31
6B/TiZXhIFHD6QYGmGdxllOBniGs8GT4P/cPPrWbH0ep2kf0PpHWUyDeiu2+R3zY
yx3Sg3FZcw2pSGzoESLUsXsoqa6e7/ME4HhnePOHMwBeipj0pHfh2Zxx84cLumkx
Nl0Pic1JCfoC0xNBUnLz0vpOOEdNusPoW9yQ/IApmJvaHog3iByFnMd2eCpZcx+i
rxswf/RoErUBA5q8ceJbwAwGLGHX8F7l1N8xmIm80QKVIb+iJckaZDlx6YS5lOO2
2wyjnjG3k/I+Ezqs3syLLwiZgFAj+MVbsCxGrYJB2XBeFj5f95UDErdM/lRqhbCa
VGzihVpNlASy/kcNp0gVDXqoqtixuPWZXhvOVusC8vkl25Iyf1WIVS8bpB6vepdd
ZycnyajY34AFlXuWszj/3FvEQmMjKvlBKpnmI+zm8K5AWSt2Cgzq4WWGtK2HLsol
QKYL3hcScLLUnyrZpX5TKivro93pprBuYKbe2hWbHeukluNMk+++VSz9YDzIWsDT
WRFlz4XmpEM0rzGx+jgo93LYaoPUqp8suvcjD5Vh7sRbVs+YioKHBYMjSH5BNc14
fvtjfnRCVPsDCZO4US4FtMoWHpsizGtkKcvpu9oTNLpWJ1ekheqnrsVZr61geXY8
mCQPU36OIvIf+wwRd1b/dFl9ubio6Ed6QKXl8eEi/4sA+HptdZMMB1bLCPtyJoEL
VMyXln7R9/Q4HroVAoplfi/uB+StcppqISj/wO5kysMjeKtcQZOK83fZpo0tgMi8
ArYJiqDJ6gissHcNgT2D9KfuJawfKHImMoE5uDLsurWWoXgWJ3sujlHocbcBQF8I
+0iv3vaJN18RNWBxKrmOxJip8Z37mRD2UZZqt5CGvZLGnNDmsjgwoYTUkNRUfMD2
1NVbtS0ITRYabXdSd4o+JXgYLgPBKomU5keJDCpgXqqBhuhaMgJgX8N9m1aC/FLm
weY8L1xoaRufNvkshXrlZ4ZJ9GvSJ4fS6YHK9lAGTZw3C5Y5xL9iqlk2FpjHVOxk
x8a+BprH6hvXQk/8/Xqe5OXwt1vAUxIsuAgJ707jk2EqZwBzP0JZtDbxpi5igeq1
ZXbOJpcTK7IPy6m5bQpLJfjz9CPkgxS69T9OEOimaMC6p7oKe0ul/efDQLLRy0qK
oDMqCygU8mueCRXhd1BwIm7io3CLL2ydcI8vqxNbzOl79Bj4da7/TcQObiEYgKO3
80p7F3zfkK61SdT0CArJiQuuMhEoBlJqFEVNwIXzKxzilStSv5oc4sf2J4K4pxFj
0dr0Uxy220u40ssukEiz9dZTF9wslg+zBvuskBxYoqURqqPVOKEfJi2fpdFbJ9VG
4G383mTK+x1OPwTlwjiiuU8R9lFjUbh4W1N9Rp7aihoQU/S4ilcEKhcftzJIJ0oi
NWOcwwrkJ9H2RTQlev2RWrT2jjTjyiRy3AtnD+XiS+peGuyvYcZc11yS9Lh3zGdi
2ak9Xny550qtIEgU8o2Y/02qkTogwfFiDcaKN+4mUNqqgI+7TduilmxHzBw3BM1s
Hyn7Xw4fUb9htMTi5p5rAVRlWyPxJKK8m9TtFIwz8dm6NfVfxIVl/9Ng1FeA6Se7
LJ5BUfjOJoqrJm7B0gfCh9FNem04FbuAc3BpWcw9VWvOayyytyyhKFcX8ShX5AN1
+6vmF/aUSlaEqlzJiQbyRAJrlYM3wmOoQq33jvA9/RvHpwEX8pV84t0EX1sOisVT
sWJ6iIKvP3gAswGHKsNcbqilfpi7yIIi9rDQ/hCOWnbyBmqOEN/BXkmdO6iDdac5
GJAYTg02TVFEQBZpjxKDUIw4F+KYiDdD8k5RzynOGtCH9jXX0jtmzsayHTCDCVNm
tTnRB2+L7S9obHEIuwP2u2KtFeInJGgMMhKxTTwC66Htbx1RKjSObawMYIZBS9XR
VkezLFMoSzsC6BMkDhxASHpmKhP//1EH+fDiYU9ftUjmrFRSRiKoPGm6IhL1xXuu
n6eUhGC+hovHYdQOxZOuQqhyC+KUdiBSHYDrR2GvdnoGiWXTM8pMvbWadNoT8KC0
gx1azJkiHo1zKmHvOBkXZJAZYjwFnXE9/TQsgB7jfuIHL/Umjx7ww0UtlziVZenz
3X5/gSnoabPbcOaSIlbGYWGO+VtM1fGOL8rnh9xrC8KfnvEDsIhakjTOQnDAFhDJ
z4oqHuDJnkb8jKHA4z98nhPoq2FGmz3ehopmwWKVAPc+RnQPm3Gg27UL8W4YzWv6
+rZQvYYiQSpqyBsWsSuS1wJ9lSAAzlTT0sWnPrthXh3oI2avz63PPhz1Fys4oWyp
DrEkhmmnu3/o54MgcfQpAGRU8w5U2yPN2sK/NPGG1EH2zaQelDwOTdWzUp0AtFrL
c+5a7bZ19/lJu5tBqGgjUooByN7C1P3kvl1IG2SVZ5CGiqxpzputhcVa59P/tQee
reCBkOpOYhNzleA1ytedS9Ui40GlORX9kgYzJSOEwZ4BP0PTuuCgMJnnTXCWrd6V
dSCuCh9n62uTjFv7xB+Eo5x8Xo4s0KoA+NTlnVPIlBHbClGCH2haXsQBNBF0/ZJv
nWo+kNDntxLVl63tTiZ0tBYH/CCUPBiW/BFI1Q5+BeKmxT134utV6xQCdr/M/yE6
WHBjvWoChND1prvVbmdmXi3VRW8v6HmTxlVTldoCm1Bd+VFAQhplGrVnFW4QZFs7
5qfiZxOH8uPGsLqpnUQOc3CmnhTXWF25frFsqMktObqVPgBcweIOv1hDw6JhT8tJ
eqxrrOMaH1Ks4bh1MOM84AhuI3a6MgcqMwL0B5yDt58F3Dpam+QZnq25S5WwHZv7
Gq3iF9vBAjmHcG3TSnnkoQrxU/otpSehuftRnhu0XA6d9OTBo+HrKEG9CumJnK0s
/6rXcjftIBmxJIBng5NScGnVIsOZO6jbuHRYgwDO3ePaUXkRsP+a8S/YyJj+0t/B
Shmi8aKIxNQy70toszirUAd2bT/jaRF4l9X9CxPJJ0eiLmR3etMLWJxMsL17/EeB
AQ8yekxw2OopU/vUSZafMmmla1Z8tguUGBZOsrUY83nk1R/8eoZtfjMiyJ9pmTtG
SU5F1mLf0ZbAjTk1gNkfL6Thsz/utx00QBNGomqF2oo2JI4H5intuZ2salaD/2Mf
ZIFRKh6m8Wr29c15LMf7b4x993JRBPMMRe5A32ymRVtTyqkpSuYYiBEzTui4dlWg
z02Mbcrp5nH28fKc+2et6o4AhSuAGfXkBQVf31ZMdGPZcFsCsqCV+Dgr6obABlbT
tU0Gm0qs43KCpUZgv9AjF95ELqH2Uo/Kxv8ljMiS8tMH3f2OpTfdATb3vixLLgM4
B99ZaXqoxNeIUJqgqaEXOASX/ysI76Ysi1ejdrpejb9Vihsdil3Odjpm0WTJAhXy
x6IKh2YHSKOHG7eWzhX32BzufJSjoaa2hzM5NSlrMkXX7ml4DKzY0aSHLbpNP685
JiHdDPorhdzTSiCxe3ATWKpFXJU3BAXWJ5yCUv0It/qNLHNFxQjQJFKJ3+WIQHFd
DK3wiXMz1Pi74sImKDVMwx0+IestAg+QY2jJeWokuo7Q/f3SnJKlnwhjJAthVy9e
UOB5vQWUHZB229jltHZB6AJWvRue47drRXF1oHIreruj8OFDMJSM5FF1PQvUvoLP
e2gemBlJ6x3cyQ0ROZoKGnnfFq/ExloDcHR2u/KZXMtZW6gTx8nU+lm4gBBjw6sv
WEFije7wO8gWP5QRITAf5FuI/25p60939p/YlXO0/8rWEIQGkrfxszd9EOsr6Tds
6nPe3WFfFCrms4TTSYCBlybuzZ2PlDw2x/6960gUpAwqz/WDeuHW1Y5NZbn0jMxj
XwnLTFWz+kisbrF4McNR/vPqBnKxxIJDRJXy69G59sD540693cTVZLWybEs8Yusp
TvtqmOzQBG7nP2ZUxRO/7d3MQ5ITIBq/oZOdUuMSEm5YSQX7h4E0o5H919dxII8T
NCm8tNBJEC1Hl9Wuy0+4Ctp/EVZesDg3J2hBzGh8IjYUGgHflIsENwDFzW8K6Oyo
xNWXNRR6i2wOzmUyaSdPi+GZl1W4gQ4ssoWPpqXJ4oXO3SW0qZbSjUOUwibqW6WL
d33NS4+1xqFbX364FGdibhO89Q+nhl8/L81dfL+r5dVLCVfJ845COfw+PUVLXhcY
oiq+w7jIxDc8hkiHe0w3cmoClCGo2ufiF/ZW0xwtNBtyS5J9mK2AaP1XpvQRAI+V
LktwR6oRULVhDTjJz+5LQi+drED/AE8gqPkxd6aUe6dUrSZBugv9irbKx7M/14BU
rL1jTuW3c3IO242C4z79/TdAeU/JIP6c0o1bRh5kW2zAdZ86iSu3gxGPzFaC4bZ6
Ly/t8Xu0KAYZGSP20kbr/mLEybkRd1q2GSGfhfXzyrxG+5tEif7UWknMa5N84wdn
/iLQloA1jcd8dthRAmVXRsCU4FEhKytTJfP7m7LVF1C7D+Y5L7cyNrMAbuZ8vvYT
VVU0JRENAvMjiQrhGoER0TR6z0g6QMHuMqWu8SsrtZOq46Gfauzl41C4REGiP68l
EIE88nT+EaW5GyIhdB3eCVyydtCWnx1Rn0B0rIKv3U2izrzGbYG0pn44tnnM41Ia
BfyIA8X+YUS8zwVq0Ir1USDkU9fhTPLczeiwxqPvzNnwv9/fm3Os6vxbjailLce6
t04qri6YMcQqZmX9COqXzdkxxN7bxG54aCespwGtjfN/NLAp0SHVw6D36FjUvFYN
ixbGf7hA+/p4BSnK60PqZCZZAL/MxNUQYnppyREIzRQHpvSub8y1JfPr9/Vs1yEz
JLa3rEdfzRYuLM8YQzD8cuIw/yNJb0Ejs0+cfpYRZCAp/z/S4SGqqRqpXKsXyJd+
zm9sy/WO2L182N4hf+ol+MkLOjoLCm5TMgzK96bsbkg/hh8kcU/84AIXebvWIRjF
lSs30nrODgtR+R8bFRBVrS/vSFGbJw4GTWenXR/sVp0EwxQU3C/Cusu1/vD8Nl2T
ZU9j9IfGZ2+HuTJxOcpwvm2tiAJowHAg4Cxp1FWxy267Ur2WrF3Q28n3mO+G4ev+
cMhnIEg7XzmkmvYU7OidOMYlrV/sWjAXuVqNJGxkQiO1pF6Y+jbYrdW2UgpkNeZV
YMJwoKqdKDg73+c+syACyKqTGedIyuMwFchhd3iZgVajn5kc7Lt+dQi/QiX+0jUH
A8uUfE9eXU5Ple/ss/MoPgSxXcsIq9QCVvmCR7pV+IZB/a60Lp7CpbFfhxnCMmfP
DjVXgeUPmJLxAPhA31SwKmszoL4UjyRRkLniDnSESOPwvcD0wASEZYMMCFQHyJNy
sqfNiLh1/n8raassadAxVkQ4897n+4oJTDAbB9eOiNOmTvMfGleca4KU1c61Gjzq
mLMJWGnal1wBSydrxAALqQqSgESB+pywTt9JQbcurKqsw31QilGityBB+XZcTCjS
1W7V6oaz9Db42xlc/Wf5EMM2++H76cyXPl77zXihFFbrDaYUmLmmuFmFWC6Z1Xfm
9uc2U7XgEu+pdFkce/OEMYo+3wgfuKZUFS6Gy9LGqEVoL/pNbWqkfnD/rzt0u4vO
u3rV44dOdTi6CgxF46KY+zqywujCUYrLmG6OwU2e9AnzWnP89qyBQapqSY9uGMhv
5pW6bNLhFfTsFbxDJgwdFq54Qye0lxUHSvcVk3QsVMgRVllcbx0hJCx/PzrgOBRu
CwngQQbaiGLIGssiNFB9o3JKoy+XCAeuRulZ6rtvTSaf6y0QsFcrQWkRaBL8A8si
5mZY1B7YppJvrvZCWnVv4jNVAAzB8hzVPiiXn7vEe2EbKbQFyn8R1k3SMyrHwz5G
oy5F4mXQ0qa8reQ3Pgszw6+72YKUmJA95PZ/XuPiFMp13bXHCsepBp8G0a2NXidH
1kj92BgvKWLMuLTT3KPgRVscPQDCywDXA5p/9m8d+AWcLWQLe/26pa6Hw/Tqq7l8
gsBkZYns3vVcqOG4jGRd+nE2j1hyeZIrfrzFt9coy59+xcJkr7x2h8Dzbgs/1+NY
YCE0hAYBIl07GHHVBDM5WgeOz23cy/yhdKLdgcKjyVcA3RGXjCIGxxNEKKWtJaIo
9rGQmiPgmPIk+2GeaDACOGTqmU9IOESZXHQNnNc/NzdxZqeAzWgo4q8lbddzgQIE
XITCnUydBTXj1pc10knhlT4s7errfSLTREEhiJefAjBkCRpcIpf4mrlYp0FKfsqc
mRovrVm5GSsngQi6l6q+JcCJH8n6r4dQEw87pxenL0otJx5cgxlZFp941SaMtcDM
L5cInWQrC3DhlK4bUwsSvKtRogMeZs4/4Mrt5JYq/0GpGUyKLYEwqJz+TFM/czsp
t1OXITwjDjYyejC3v/kbiO+tTq12LXSaiI1qcid4cDVQB7slvD/aOLrbh1WPX/Cr
ec7QhJKmwkdpqlW0TTk3kkBuOeix8NT96SW6MNiR2dgF7ykqz9XbY60DWeFoPEhg
F2XFRLaY6NoQ9jEgReH4WR7BNblXUrxLLcxUZ++ic5zKp1sbpF8KZxUK2yKM+gE5
KY/+V5I9FXRJ4yW/j+F3QdOwnPymcDxIcYVrQMqEsUtQtKamBklktjU/0jd86UCN
EaS0+owB+Eq0SaDJM4fJk6c9LopBzQ5YGYEbynJ2JAFfNASU399k6n7MZ1ao9hxL
dNvhA01Qaiu/ZlVEDFi+v9GMdQ/Ok+TdcO7dVeUlRIqwfTjE9A+Y4S9ZogfMiBrV
Vq8y2QSWtCuXpLzq80KvdfYR6Tm5OkVxUnpwuEv79wJQPr3e7Yp+fvq6Uym/g94w
PZFd1RxTdYDoWVv5KRQNzI0qWP3U34h8X/UxnZeko3yTKBSftg3gQJPxE6T4b3/m
KH4KPHeL9JGY9kN1bC/09SgumSNaG5v9LpQSzGgJn80S1ZrcLB1dWj2PtP+wBPtv
iPJGJOR5v85SWmvLsfPfTNIuu9HD9ZlxruGaC8RX/PeRZncGiwhHlXOHy8rdhe1C
wjx+uFRdlKK7zdsjxh+D7+e6IaJ9/0lDEeaGo15mwmn0gy9ucGAzh4CXJRxPGs/s
CPdf89ap11W9ooNi2eZPOSu+u52fcMzMVBMUXGRKQDaXnDJl9kwM91OR8IfwPPSy
BU6OfJK1znpVXKXcJVyyzshyuOBe5+HbVWTtbl27yGfTqoy2yx3wYXeYAU4n6IJ8
LcHM5R1X7DjxuzjrG+TeT1drYnHF3GUYzZMvwmQDHTsWeRR8cqEHuR3ULEifa8xO
mxH5w8EasG0Qc/WiVHyVzkgbrFDCZamGDmJBvqKV0awlNXjwTkykNzy6NzIrRRRb
OujCPQexmvaphgz43kH/FrhAqmlLaboWdvIbnCsZucEZz01KH4xBEGrBSx2J3M+j
TnQnO/FIf1m5FnfRxNpAKt/tS9GXCfAueld1UGwQm1enh4EAKesq7V1cBieCDIuc
qT3ZLZQtWtw62ZpOnxdkqzSk2KHvrvWU0/hArZwFQMEs/Yj9MdUmMG4WufbZTtki
rfPadjQILXS8J9tS4WUcdN+zOdTMMW7OxaUb7ebs0B9kHNj3matj5NAghfrNn2co
7WF2nCD2s6dfX2ZYcNARJeybwX3FeOzU47yUr5yf0lVmvStbEmurHxtQ63dvR7Qj
GRvedgj3c0ixIaQUlzrfesNelUvqrpiTHbuBGErebfb2pv0YjtBO8FiOAN0uxeG3
pT7YT1OWpAJRg1w16shfD5FNARVKpPTDa4UzkajVaCR/kvY3f1RmdHyNHjxiwggg
5YO3yi3gah5cpyfGS2Mn84MsztireQ8GEYTGiEJeFcMJBs9J7fcaCP9PSsvUNBu5
u7Qrfpt/hIy/zITmeDnaEH0rIfYhJ3+hOSkr3J6QJnNSRiPlDTZY71MSGt5WO256
qU6egxA0aic5debkwZP7mJPkYudhmXP3KsXpJrBMq4cggnP8QO8VauN3M1UQ0lfE
e89a0fGOlcO3jThX/KzeBzUxz10X50nKBeGFIkiLajkfgoBS6TBm5jz5jD2Ymin6
Zm70SbzadnXYoitMH4hhurVLQlcoUduuAedvck8miQEkNs4XT44hTm1smFQxWfS2
RzIXBu03DEpi2R7J/VuI9VrE9Pw1/6+VFaC6V0b+/m6agGfYt/Yx7RdICa2kobas
7jHv/Xy+8pNnQSVHT6G5dMJp0owKtzIMqlYj3pZ0BZ2rG/rNbEpIJDlMRb7rR4iy
NcbqaJuKh/FiGjxDL53PFzhEBgy51SxaSuOV9+JVeL7puxZIIXRHULq8ASJWjmI1
KYwSLJcFREfG6abZg1+LyLmJg99L/2fAAZaUeFehPxR2jqjzvWcIOmp1+EAPjPVX
mF0N4nqQ4oSWKSopsY9WP9vRoqPHRBpd0+9JDiEdOTJGcia1yjCjBVc61oMIQ0NH
MIVzlnRLMMiZhkewcrtD0btdB6srkpynpGmSf1lAe8anzbHDY5FnFn6pdZcNmRum
VX9sjylhatSM60OzqT816gGpbShD2NQ5iqXrKHvzB5tRS1FieHJKpN01X9FShCxp
nN+9B/k0J6VhKkzJjmFU0io1aKLQ4k8ceW7q6IGznZYwcMPde7Ia2VakQEpc7MZS
8nPTBdodWa5adw3E2/hCHqOUJXgMc6Ll5pJsEXQS+X0lAloy6BDYtBpggLshYIIX
vbVrK3CCBXWuR34o6/3Dgw9dVCo22IxRfQiGfcm524AugcXWMFfBtfZuV3y0dI8V
q29Ue36/Iw70csdliuB3qF1ELDXZYOAe6RQ/IoJVTJ+9PFHY1u5gxQdFjXBCxxVl
Y70MJ5JEsYCO07ODB29jmviq7ivJ53AfwP9DmJpdykzl6gz0za3Cza6P9QS6Z5Ih
Bq6rCA3W8PhTQHUYo3qMExJnTe0OdZPgfUx/7ub3WyQQdY/akRinqMxxFA8a0wrr
SkSPCAIsCl7LBSKphHe2Vn1v0MHyirLw8ZxiGxJP/GHsPC1+UXcA5jsmY8+tTBw+
mGbqAJu/CsA2oFCW00gWac6TkboHHjYim8mEhwB+EUMmNEF2Cse/ukkYvOXtNRSt
Mo6CO4WAJzFXNQYcwplICItrWc0vhsbDlVfyD5m0QEXSUIKgEehBdJDro028IHzB
e3rbgTlpypkdtmNOt7MR0bPv2kIwUeLSNJ9Hp/SfHqS5JA+IVKnRyWLoLMRIVhIE
wGYyMQJdii46IyHMGwpDZV1eXadIojMD57RWxE1zn8D+u7JIxlSyp4/PcidMcKHi
qBDYTHxEMsA35KhmYxi9iJwgU9IiqQ5PFNAeYnnupAvD2FHslEhog3qQosLjYoTU
xDUqLcIJ7jQ89dyG+7ezbTtk8KcaoDYTkTu64rFlLb8DqkJbkXUTs7QNkKKnNb6j
BfpGsP0VjnK7/BJJ9QvQi6QvOolfjZr2BOUJEPLNnKagllNiAodrb8Dfy5Dey1Gf
IYrri9lxkSOzX1p8Y3PS5Beri7IssbBxi34VMv7QaztynjBYLvfLLQyV4T+R0ts7
rt4uJH7cLTrAbxZY/soJ+qcbARKcX9y2e6j6eUrSeXRnE043P0tGiejdedK2r9Q5
QJPstrY99rvcz0YMPCX1KFhasr6K9LlJQxathXqyJCwysNs/ue+OgQDOxOqElyQb
gbCfKjcsBV9MsnVUw4m8KYFaOdpf1FEEuQAHh6Po+JSUXYebvONBOapBw0PS2CuA
JppsE1Yp4yb6N+tQr8Ces6UM9Ypq6Iv7D7LR498ff2HTAVKbFSs1Q/E44QNJ44wj
y8xygdo6dIDjJ9jRhCHY2rCTFxU9o//uMBFiWQEgbeXAuwyRsXaqB7VrStevQIDF
yjFS8uM0Lrt4ixZmu1UU3iOEJqcCv/7TO3zb23Pg3qUK2kb1vfDVpLjdmLZ3wwXX
2eSPY5Mco1+kG5UCiv8P6Z8ioLkg98fGo8rApCXpCm4eviLXAZJ34kyLgJLgLKN1
mCh+t4uBVo0BfhnL9c2e2bZmHdjvaQaTr2dczCNzqZo5wTwxDMKvnDQmiWZbtMT0
Ea+WA3hTHCly8tORYQYx4MWVfiRN7g1BVF90R7vWTahci0mKwbu3aaEBmST9vDq1
iJsP4xR5k9TdSMGB0uqJummgw9GaHnvyVXFbaPipwqyTr0bLOSRsksoHlR+CMyfE
8aPZTrN9hxnRfNn39+lLLT4lFRIUHJRUoZeJU1zpGkjTvaNNclpSTW5YSJ01SQBi
KJxDS3P6sUDRgqFzK1NcFOPJolGBfFwt+Tw+iBupR7dR5PNkrjzRhV5LUjBvyC/w
rNqPWYAXHvJElwtK36qSIl8Htdxo+gH6oeuxsXlFZ4OCKDNUEItNIvNMSoiew75d
VsuKL3fEa38wt6V+J5t7aO9tmheKeza0ZKhBw+Kza/EG2SC8BLS/1WyJs/j+CQE6
wRPiBidd5CLB7fKGeHMdlkhhMcQA46U/G2WrQE+WbdpAKSGbYIoHHdFFJlfDLbJG
YKLWkLeA+oHjAMhG+BLqesSBm6qcB8eJOd5Oa66Ewbm5tOTesMauHPwcVQFYJtKB
O6larWckrUF3b3gzUZ3SozZ4jkKlI0wxPs8B22SgdLAeKir0/PJ+B0DDZuHVfcKq
V6DAvfBskIx77wy4wTlvnXLyOeu/zXy341YweLeRFT1syG/rJu4lLqDoWMuoMeRX
/QXbMYw1a0qBcpSfAqn8yfLfyb5qTtm7EEP504MZ55UZhpxNxlPnzSh9Ddj7Ny4L
d241gUyR6KXJuBNZq6ZIO2YlCQgfS7VyC2Rf6hdrREDdLrjIgAdFufhxO5roEP+9
dErIpxp/a5ZDgdgwMWzaZj8rfVmyi0Yjuw56MPEoew4+EVyfXvOFjNVEe98n8Ox0
HpcNIdL3Uzac+GxUBjfjTZ56ZQf47ykXyRygpo8ZyN3iAqnXHMfZxirAUjafCrYw
3TPjSAzhwRp9DiPn+Ex7DZFQWYxkxzZIft5KWxMRfL/OpqNGqXJAtH7WFEoVMghe
eozoIRO89oAsLWJq5jvYX/5Hc9l3p3k8UfKuedjb7AphOMAhYcuhGPxFHF/SALjk
jtQ4/lKEDMRaOXcKMzcAEgEZf++xPvaasKVAseKF1V1MfpuvcbD2+XcD9DJIb19L
EgyOlptRYGegn6UbocIM0Eb3HP4rsw8h+sqdeo4BolDtOiGbmRIAMkEaifjarYg6
f9DjdDIwFaA9W7j9GBBRLFsVJzu1VBZKrjzGeqeIaxbMw1a98g13qeYSrzx0cqNN
71ZPZkGIqnQs6L8ww0a1jhIPycFnis6VFU06PVwFInJnJE274069GG+xBPe5OTS9
am8vhmsAjRYERLtJ4F0pnde8a0fMkAwfbGOcrThljwoa9HTD/OvQjgn0l3axKkcw
BfU/+gcahAa1U1h3Fy3Lvk0SaGL+VuEfoEpD3HQ9OxBBJeomtdY7PBMjEZYxd/o9
ZYfrImIqfeujmTNVztHvIm+1qFoLxW9ZHLirI5upzzmD/5wpucYZ4x19wbT1fNMY
LnNJOhUjrEb+bzyEoWJg54xccbjWVW+rsdfI5iz27AvILnMHgNIAVDh5AE7X+RxM
aOxWhi0GL1W8SJ/0duxUn6kHDljW4zt49nMsfhmOrD2LJ1YbJcyINYp0Y1OYj9gJ
2AKH7JwrInHfcGDweIGACgcba3A+yGg9IqCPMqxuVfcQFJdvNJWkGhPK5ayzOci0
++xYwybe2CEP8UIqO5waV9uqQYbo8TvnPds1vnz+zx4kaLnh0T2aHiPdvop2ElUN
u2uawwtW3Tz6XXLEe54MkKHT8bwkjRa0rq01V7muo4jT2R3N5v8nEE8LOXirMKkw
6g7666e+J+4tOjwFknQTZkRkBqXKUdnl7SpeHLNji0T90L5MJov1B9/qQ1LlAUR3
qCE1C/MKRD2t8RQUDxRU9e2DTX97mAXI9CbQCoIjRsP6LTgrqMDkj7HgVRQCHMZC
kHEK3NUyX1Djkjg8kpuSxu5+KF96NjC4dW0/03RFhgwDf5nX3xa7j4yGbXfXP9/2
IYfmqDgwLnbmDGdVoX0CpH+EW0qLHMo4HAOCL/44CS+jw9Yy+a/F/sRiZp5n/0Qp
dZ1m99U9xLsnOK68CiVyaqVwwpofddSPXOTY4ogwJkS5p2/ovDTJgQ7dvo602RNY
ix/Dow1KuCXUogui4wMEIvxBKRJzyEvY9t/4w4f3iZFZpaAeqTsa5v+TeY0aT2g/
W7Ri4Ue5iZNd4UPROkz0bEpbFSh8JCU1te8EU3JQ/WyCuleQaaUCayTNfhfr5LMU
MSBH/3L9Hx6U7/CCv5Z9NSZKN+D7FonYw6OAYqKcMSfREOp4zIoMflQTMrtODFJz
mzXo4ZETn3LdyJL3Kc0pj0wDgb0y+UAwO0pXsFk4fgHI4PkD6oMK9vZqE/kimA1k
sgKjWQ7n+Gw0VW2Lki+2+PVYibUsQi2ap2JXMwWmeEUCKDbpO7QfWiT34jjXOKAc
2dJV8oxOkqqHAvTnUiNGUuDjItpR5qlNAEj4tKemPa7o+DzkujbFjdOfr2pKopIv
OqBicyMmJU9bIn8AEq1o+/XZmOecysXLZuHmN0MreGyuxAQKqnD7EIZKOX335ZF8
u5yC2vGZ7JWC+52jYVZC69L+WH7q0NJwaOEz3YDn44bkYgj2Jm/WhPQErkLnfiIH
Iz3CyvAsxAhM6o/F9lftfanPUjjych050igaS0yEGBugwTue2JnSJ+j0BZHlFnRV
rw5oKL/v6QqLDn6ezqTk8qjfHO8lxIglwW3rzbeohWlpMx5jSNAVXdVtS0V3LYnD
6S12TrWChXEiledVCKWsphKWFDMzv77OmcOFBayK1454q9FT+MrCx5w9TyE8UxoP
6+tCamw2LGFuVbaMPGyR0ZWzSroJW75k5oNaKXzl/xiZtTrNr72v8xHHjgmPE6cM
Al7IRSu2x2EejIRAk7XIStqFONDSwDkR1FuZZKSjM/CAd1v4agBYw8E5ku84XZb1
qavLwEHUSVlMWHCDQ9iNisQttw0KyM/CDsrD+4keMT7s2S1tZ0dTXSSBDFh2psuX
6cYDVfflfOblx4yUrtUFbP8svon7t2lE+NujYG7fdvCmUAj9gtZdf1l3bRca81uZ
LK2dSYvRYVkg+Q1SPZNLCyOtmpZ6e8nNaV8G3PAapd9OIkfHRSWt+q7Z/u7llRj7
5ncDSzQG9FdXwbFomZLeZxpPmsOtc9pa6lreue0ERXxwW+rec4IKKl113MuZfu03
jb5drj/J9cn4DGsf5XX3hdPIhNJfCJt8L/V+c1b7r5QN/jy+eRkTor+4lwFcxfEk
qjSuVG/mS4KyW9nerjtI8ZYG9Q56rJ5FVaQQ+n7b/PWisMO21NZc88Hn7sV1HINo
j8bzMiZ+M6NVmFHEp+AqitO+c/2XMUY3JEh9azi+5bz6BSNUIaGBAzU2a03b0WIL
ayiqedOuNYy9rvQJAxorQG0UZCWv8CC2VrrCGxRcKZLoG6s7Le352VAK4LHABYgT
/uju7sLn3REKU3oUaU7eu4YNYJ2LXwkIEVtXyOXlfY5+A1tW9SY4TmUeRRjxcSvq
JDwcgbH7PMXfCNfgfp/GT0H5GOISG8cEVigFD52EYy1PALdltGCrgBAV+gLrg30u
z2Bgxv2L6mYldonA9f6nYNZsqiGAias8oNkfkA67tvvH/+NIfdx+mukBEwl9WYFW
HzX9s4DnD3mKCP9WSb4gF6szsOAogJbhs4A9aJtQBJOrIH+VoNVkLk/Pt2o//0ZM
zRanI+yUIXmU0gaK9p5ZmfEHm4O7i3z4Gc1hXo0XmmvkXDgKN7GXyjtz6SV8ZoDK
czp/7xKiSHrtg0A3iL8RCaI5cJISWRiSpBUF4S0L5Of3nWvBUfPAjl/sxPTqG1cF
i5yHjqhCho9hU94/lExnikUCCtG8H5EgX4r9FFwZqePoQO7WElD9ion2hD72osnU
j2cDusgBRE9Xteu9VrbKLxJlF8yCV9bjKMLSg5Kq59xepnloPMsvUp3txUaNdn6F
vYlpiLHnvVsUn56JopNrtHRT8B0j54UhxT3w7Kz2Z/Jdc7eXeJqEIML0bpZrmOW4
lqcRN0YYw6wJ/JTm5/OCK0KoByFzKWFcl1gftE+8ApQhLBIPVNp/Yc2/Y8N1pqi1
eJv738SIfrlVpVc1wEwqFHRv6ihFJU5LH4h9Vuiz7HZcNnLGHmTBmcjlfRtika7f
CPclpIrmsfNy00NlgLFHp53KOVHS5OlKtagCjz6iebjEDOqQ0bkcWui3+yXRlcd4
gVFgTmrzL7LgygThexxSbCljQXlNoMJ75fYm8e+TnejGEMjZTK8p8TfodQfngPDw
BKezD1pz5rZV7+n1203Mz8CBMaM1RgCnvjVl7GKpJiO9Dh7xL33Aarb9XUKroWkR
Lhqs6CODnQ3dp+K/2vpmPKbD/zq19LOxd1oAO5sMqXjEGloUPd3aOBqwxing4rYH
hjlpkJrxDkL6cAYptBZ1PfzEWRfAXgFy4T7RIoQTjxgMuIrom4vKYEkgKPSj+YAn
0A8niTW+IHaF8FAvNBlWpvc5Xh+2e919p9WnjDVpogF0ufftnZhYuVZYjjRG79DB
0oe5hsYhtYxXLeXRzZKjiNZmFZNkC2EjXruzB9z80LspIL4htrltmUSWwEaXmRnZ
mNXfLGs5w+HWDX8cvHeqrP/qhZ4h0eI1pNTexgWoJb7JEBOuosBHVL7A5vGUyvyu
q8wySc7RjJQ3d6Lm4NaiGBR4ShU3DhslUteXsr6BomzwSC1ad5ckpi2UHhxa/TXO
OXIEfpr8oUNAK2Zg+0QspojWvJAWiQ00QbQDlKBtr9EPKepjCS6s1xQdxSXvDmxs
6t+okmtWRR5I4cEQzeCnC8LmYltr60d1hsYlhBHN5X7XqEgBoYnfFdpCB3RqI/Jx
wbhyP9aS68+FH6ZYGo8IzkEGOJaSXFl9vD+pUkwPmdXPkTLnWYNngWOqYJsaZiVY
kw5CGxX/pm0kfJdAuqvGzQ==
`protect END_PROTECTED
