`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfygm+SYius6Id6Pnuc1w+Du1oE0bJ6dIR/lSV1OJOgv+XyuQNERAjXO3oS67cYE
gLCyt3IQ0h6kSpe8AyRt2mnYln0SrIYJ7NZsWfkxuFm1bEbXoBhhdzw/bsPeybAp
ohsN90X417DUWLikmDn7cG2NDUqdw+IhKuKJ0FOa1/1NRith92dKzK9WXEl1c4gH
tyqKaqAFr56E1VwCKpX0+HGUGhImZ/AHZ+wAfsddZttjqGLGn8aXdBpMIK5rc0ha
LRSGqrptUtHZE+KwJvW0T+S/Qxcaprq3P8+5BiKBv7ivH0CTMouN6OA6fuKsK7Iu
c/727MChkv6WNeQW1W8vBgmNu6msHHbyVLN66Uanm7g4U4CuKAcVFcXFAoB5Xhnq
dZTVDwp6mJOZcUldOXpfICaSXgV7uZGdW6xO5JRU0rNYnTnyBbyWRbIyUHffDGny
CbJ7YL8/358DTYrDMpryaG0F0l8Idlx748uOFyACiAMyoKVV4neutR+sOuPz5uEB
N4pssEggGtyN1jU8HMewKBNxKr/rtyS3wYk25FyxqZmt9r2FV4I5CHEeP1V0OPJg
2VhqBOMf9iwX9qUymSc6LDjNUGD06llDiNpP/0nBulhAqmTCnG/xqziPWJpim2vZ
yMoejjMLCsGHdGxjHW4fBpF4A8QfycX/x55N7TWBdtf+RbM8//gOTGY3ByI167N/
TBDrk56G06a52w/y4eQGAMfWOxOPT7dh9mzeYMTaTUxSF+K2lUdXaaNm0i/0FO8t
+LdII5PAu9k3ISSWu+Oom7OzqTSZkcs2G+kiB2FMlYu9yHJSsbfNUc2OQ1evZ7Z0
EoLMfJbeIT4dvD25So/XOZdT3tR9ecYzd9+FmeSGJ/2m8UYrIe4JtTbEdyvLThdD
yPZcKQCJqreKMoFN5rtPLkXWwTR8KKnsTvBHHLooKvsy+1JXR6AQM/fi1j7G2CzD
UjtwbCt2ssbac6PgnBTKdpgc2QFN3HqY/r4NANjs5FxHmn++UOdoaWJGaiYPOM7f
mt0Bna2+qYqclrESeib6qfveGgl495lq8yMrHsBNg8K5x+ZPvkEfWpIAC+wpHo+u
MFas9hkRY4IGiMhmZIVsTriArnVPR6H96yo8SKNiJZrQaIkODAysWJS7niKmT35z
7y7bEvNrHuuxwhTNDJxXWz5zQ6KX/uuza48zU9RMmxQ/hse3P5xx7VWwzLuzzYjG
Y+SdfbtSgH82v4Lrwd3XBJEfkqV7fWnV53Uqp2WHz0fshQo7Mz2TRacAGTbzX2YJ
R/IVQw3jUfCepF3oDPxe4L2OrHtdRVnZOSwIXUXYt5bvyKL4PxerO7abXDxuvVMW
QU2gY2/DxGcOT+b0N1VULroztbM2x17VR1f3rczfuMbNQ7Eu1O74KQiJ45+0Gi+r
aQuoI4bf68Lk/6o2iGVtANBI8BPOY9urkyjwOafnGyUmIfAZu4e8Y1xmKrYmLYdw
T/nZ4lvtWNxlcKbaEXl2Gzk0XCnWhsUX/s7fpoHTckPAgFQjg/rlyhHmsPzc0n3E
46DflaNSLxIc9b2mufgHgQSGwy4SZgGamZmjhNsyTJDATPAHawHM95lNpBEr1vUH
TP3QTgRWLOiMPIfUhTdyel3hpKG4LmwLqWk7dX2xVGwDIsN8Wt+ZhAJJrfG2pyME
FO0tuwk0ScJ+iMBIqLDtxahGcSnUPt6oVzTG7qsctY1rA3CNetjf475rXvgio54K
IIaCJW0Vth+FQsBpeUvseBgZ8zWwhmD1dGdaOt8xWog7IzQx7vHiDkzojLh0lzhE
DE/+AZseLeAhctNZASFYyn/geJS6FHDuHLjnXRK7ndQFe6z3Z4BctjwDL73SIvSB
+dnDBdAhWPNVlN65sGRmuFcc9MZ288MsVxsRbXtSK6e4/mrRRt/idjhK1iy8TbOI
pS/E2nrRggKumrzIw4DkaD9lzCwymXgF3BkxnB5/AqQ+EgBhIMkr4x8uvPFxubFC
w4MYck271EeM+HILPSzBJrZXTGk4ZDrx5sfTKEoLNCdB+p8svtmfvkpp7jJ4kLOg
fRxBIsquk9UDicpWRlIxqJIiEDXhYoNflaUAxTNwfpMmBpcKwb65wVAPMKHAy6xZ
cq4CCelBwHS1o/GJgX1xHy4GAkD86h8OJEfeqJj38rh6GvKNb3GvSERxdPTKtpx1
XoF7bkOpsxmYvyM3Etjv69ijuS1wU+wMUkO5YqpG9w9/BHuZG6RnvVTZkpe6b5s8
6p58e86j1Z/d1T7Plt3hY7eDwZ+TjrPCQaMdKsH1GcIe7RYPFVKLGG0hT7MDJyg5
zbxWIHzqykhNGn81GFwuPKyeW6oNzP0sIHrGilEODdAjem2yZb3Xbf38KYcklxJR
e1biaBDTE9lvlPwDFabaWpKDUCyHvVG+Mmsu+jtk+e3B1Mp5YbK9St5QS9PF9t0D
338wz4gtZAI/VJl3BO3p7P9AMW7BjNv8eitwgexgPXM+QUZqErYU8+0XbwGnsHL3
8gXo+u/jrLY0A8OatZn/t27+6FjG1170/aTK8E3eUPC2QIMNpxa5n3BMmIoM/L0f
7LhRcusyiTH2DgSPTGhsRiygQq2ldYR/8NP0XHA+gOB6E3HqSZf9gzzEOYh1gu1h
R5Mn7O+/ptAmBrC8E1GSGH0vfKspuPs8Ciz34TbOkUgg6ldYNh7yjcnXOe9LnVw3
UmxCINth2MsYHxi8R5z89xYCkKvKlndfgyofHtCFvesRKzZbb5cEvAbHTol0qtR+
3ICRggO3zs3f0bDn2qnrnV33PedjaL9GXfkVkcRCsrhsO7u5280gJEGgsyKDkHcL
CrxU0GlTEBJpTOqgARcIfrZG3EU3SFMnliVLJsrjn0lj51pixhd8zWvvhUmO6bOo
J0Thpd91LXVqgh8UPjMftvHvC5N75FKeAMmwJuTK7oq8smTn4IPwe+H3StXoW0ev
GiQu/cZs65eOLiSLfoBiZ82Jm2lCfyLJefIRx13u/uMeWADUDIozlWvpjSzLLImG
TA9A5yG6a0fUvtEyh0VqYyZpv8nblnvNXT+K9GqQkTvPTWBxkSlnqGOnnXxbMA84
QC2RDEWFGMu95L9vYg4Xj+n9RAubiWGwCBKqfTqJmHhxQGr7SzH7j1zczVDDLvt+
n/dPo2G4PLjmC5FbqfKE2393gHrT6LDenR0puFTkQ8vyCtHTN2ySFZKdny9fW0r7
EYzLlRj0GZKBhttkYmELBlFrsYiYMdleKKx2uKtXNhOaoZ3diq27a0njm0Ql4CfX
I0TAt/Z+1VbAO4x1wACk+kFTS4mxVuOzY2np3/uyKy/Nyqvk5MweYRqwtm5kpzyT
yEFL92XE1zk4JYwGY9IIXkTO4pOAc4R9T2NBRjoGtqIG3GcaAInGoe3xSv1gC9Qh
6ArVf0Kk7aD3GQN1KjOQ0MgDexnmWY43qomxN736yUEwZjiKHlX0fBO/X5gFoZBx
VuxvDCGetiTZfoWghHuq1UZLD8RS8H48rx7ZNLOsfC7Lq1j2WvFWMfH1gD2IkCUF
qnplfTTiGY+bPivg8VyyNUcbpvA8Itt+jWsFvC9OtzIZr8lhW4H9UPAh5vqZQbxd
84gRRM3JR2t33RQyVMML06PI5vqKxC0ohPF5PXlCo5EYlmnNc2b/ypDJiMTPHQlO
tGwmKJcOOvYpOdugBarCOVnBgf1QgsyuTDJ2iS/aTK0W2ZCnZtO4UTXnTLgB7VuH
2g3pkQ3k1HEFKmmG6nHug1dSkY9/4uHxYqjgZyjYR9JC5bvZs7s8y2RJgpa7oeln
XPoZGzfeC3IMtfyNb+ufNjQaGVVpxfC5GuuXu2HO9AKb/attestg07cbudoDYaMP
bqr/ZRdp0D1S9IxZu5NM8WpbAipnr1PZ4fZt/Cbu3qOuY4u8vL+7eXyIFRWWjYbH
mVMQIAWMGpwOvXapLGBf4afSUJ4S2QJX9gKFA0ci33w8+sxBQkld8PkFSB0BjbX1
wjTc80/R7HC3E6RF/jctPzNtjck3SB4GeHeHZ4LL2+Nnz0z3W7b77qe7CKeghkOd
sDmS1kLqTir2ebKcb/QlM0nT6vxvZKfdjihIIjZ1QVjwdtbqSCneFPZlR7PDA3hB
cRYXRpAotenziCV0kDHuXpAjOmYTf1yr8eFd6A7lYxOrXrW1KRQeOnwQTjCPLsKk
s/AXDqzA44Kt7UKb9eX4K8GjP9kX3pZ4fnUldMZsPoWz7YdJxKJ04AvpOr6LywL4
or9iIdvdrFYmlTWA1rU62qRLJc0BnCFASjfIpYKNmrqQT0dIKZQZ7hHWhqOnnPU8
7wEOC8fT5dKLdVApzWHakNVz5GhRgnwm0xGvGSxmAw1p6Rf//sEHbqsPZWWaLzQE
Uq0LGj5pLTF+tuejAdauIpB93eszkDRDncVMFfdRzhP81ilJurgEdcbxSuRV0hVH
CN7R+3AM7pqf/hvKu5Xp7V6RyLLY0h4Bla25abPWnnTM5qcviPCH5l5YN4G5GnKJ
sND0SYa5joxGsohJ0SR3ED6Rck63sD5zvPKJZTpCv1tRbfUqitH8B7oStzT516pA
Ldql+k68FjyHmfoLilyPCZcwf7JGVkMLbfm4tcoGH4E=
`protect END_PROTECTED
