`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FwCXXxXH6Xav+X9r+MUD6dC/eQam48XjZwHznV8GE2GH+Zl1DLBjk0qgq29QsLnS
7UKhJASQAOU4kBzhB2gLugoqfihqq9HO7Yvh8JljJiIQCekXzKGPWXQXdxuXBvyw
/cjJqLwB1136qasoyBRF2tKwmkwoB/AVV2kXtYgXdMOdZljfXIFACSp8WEfIIB9J
fOeSCAtrXtd/W5Sd5Z1y6jIOGPi02p4yxV3ds80OtaVPUX2Y/XFbdOx/cTyvO49l
CuVaDJWwBr4+BcA2E5zMfVFRNYU26LOggjw4Jx3zTxzVulf/6RQOXTAzs2W+B6gj
RNrAPZbCFxXjiVarrHiEVzeTlV7XyNyx6FlgSeCwXWzsIiYIClMjpy9cNoHA/NtY
wleMXJEggljJ5EY8Spa4pOwG3Tzdz9Pgzy3jMm2oAE6k6zRfDl5zaFuxkBh+beMy
zzor4dd5VJ1SOoR6rmixuJxfoohsdFs9U3pFOWGxxfZKvXKr9cqU6QxsSPLcdPXy
xVLFMBw0HaYmy336PdJ1TpKzgsahg50LpHmMiCOY5Ky/FdseeNy81Mz5zXvB28Yt
bDlWXVPITC+RCCWoGyJh0Nb+Kfu4jwtGmG4QiQPx1hm88rm4MGtwqWGYHUAouLtQ
nLoJ6+mTX6/9sIhhL4yanLOcK7jV/n2b+QFzcpiPnUiRKQBs3JkvRDmLk/iryWWO
p1VFSVd8sA0N/tRicWrStzglFA7cgpOdtYGqhL7fXE+/JOIORZ6WWiGCDvCnFjSi
l7nGN1A7XjONe1CrZgH5jtM2izBrixULyFzc9xhmwUxY9cqdcY8E6pca3oeHQNlV
ghgKJxP38nKRueZPrDY1DQl6xVGmFZCDRI13A3+zPGzetaqMPDyuCNl9RiYDhitI
ZivYO5SAFiEkgddTryhx+J41zO0iIx+Jn1U7AvKBoh6Znx1F+DE49RbHTAhOBpKk
2f+24t5060RY3wVDeJ88KvRTSKjurzsyL54qtF0ZBnqPubvcaWrK6/X07HLyp783
Fw6Z2N6gmbTfWasIA0kZONwbd/HWMXwg2EulhhlkFuJOsda+ix6NU3eD2RwlRk+w
thDcAslPS4Q+FThrC06zCbCS0uY4VeBPUW8NFWj9hrufSloLEXy/MLuefmt74GRy
uxcTaP/kMavTqWjkSUVc1YZb8XdXeXmqkCGhnSmA11XwBNUiDRize+bjCv9Ol7b2
J6N6BrqnZXs+j4cmrS6UTMft0L1Xi+JqdeHT1DcyhkjkAn9FFwlIJtnuGCYLfz1P
ndUUm78mPgiCkB/Ik5G0GvpchwUnWCZcfB84rCqrN04ewf0nSeVIzZSb/BdbMFV3
W8djvADxFrhUpsssmOhhCbzVn3Q1sASyn5byEd9piJ8oZiX8a0HWzIbfisjipypd
KJOPAAWEa5lEbGSvM2p8V0dGCCiEkgywTw6bWjesj72pScS/Ujnk2WBiS2LC4Pjs
mefh18sWVlTPem9mhbY5MLfThH1Vr6+Mvlqajope01vf8INeENPeyV5wv1cEyISI
0iWAbfN28AywpWFaUqzSM3gE12hGnlbSqWKPHYGOERRjmfEnLojTwg1nESZP3e6l
NbcvrTVCTsmVw1clD21O5Hc9IgqvrYNEyGNfqFDhYtGP7otBmSntEyT2UchnFWt+
2jDBcnaOCDIpgScUwCPCJ45YHr/T6o9XjX84ySnLQI+KNOeMDXPeUmN3oUDY4PGD
I2rFpGVZYYCxSPaKNQ3727W8VUUn8YtZuwDmFoOJU2QMRS6neQdU4ekan6mKEtOM
xJHI0f/nwiG/R03p1T3yDHAhSYxyyAQyhc0MD4f0ObiGZVD9p3P9T1IyNSnc97Ka
0ek+j/3uBmVqnlEooBHrErrSl4zOapXQOrwKmKhKM7DXjVpzziNE83K7K19p2+Zp
93F+pqWBABGkK7RW/aECTnY5K+Z38x0fzvt5TBpjvcRQSmlrbfjvIAm7X3LEjBmq
1qeayFf/Eq7KtljI8SqhpCOYuLnk4uhg16Tav5Rvz6SptQCqX9Z+jUV29si8+jNL
D9DKLLhVeAYyHqViJZUX7X/eDML24TeTPSz3ntnEuElpXrbEXUoPhrhHiaJnb4Et
faBg98TRZdNfOL7YCA+XSK04NrO5STcjrdh7Dvzuv1Q37gXKOtkAX86TkRiw1GAV
NgZVPbgNzhPcgcACeRkpvenuFKRdtA/CdXxxUL5CB3nvnaQxPbGndWpsr0xTvH+Y
ikH6jGLomDNslSBiPFHgnz5/PQDXTbvnl/Wdw5jq1Hdjd/NoN9lnmg0fbwYJ79iR
xJzQlbrACrF8/YsAv3jz8jGz1UfFP5BiUvKzvy/X3bifLGrDTe9PNEaHr9BpFCCf
R8YX+03xOKtaPlyeq6p+ImEAVRLuGVfFOAxaBbP9Jvh8ARt6i+L0chcQ0VncBBua
AhsywwuatLTymRlGyvDo1Gjve/pdbZbIE2Uu6BqYOWBg0iASrm17XHLWGm2o+Gos
BLV7ufCGvlldWPqQ4Nxx8Vt6H02+ARQ5Uahe/SwVPNRv6B4Ubsr85vopnbny6n/U
xkpmRZdhqerCW+vzlZ7Gf3shUUhPjS8ytPleNK/LlT8/Uv6tPv7+so7R3nuwpdZ7
rFrgTTJtVMsCcP9q6bkqKDrkszmIdj4HzD5a7F47Y51RojTbn24kdvfgyTj2aYGe
Wr2vcW7HdiHFuE7BTdnKH+GCr0HkHcukj1QaYMo9MqjJ4TjwQ/E3VUxTT4wcOBjI
Uu58iTLMO9LAskezTPxozw==
`protect END_PROTECTED
