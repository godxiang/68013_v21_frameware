`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wW5RNqna5Lc8GTahSmlhmtSqss+yntG3tWj5KNgLs0N3kK8mAOJFrQ7K+zkWaFgV
Itc0OQGFwmeq+fN0JaysLGoExPrCVlWnaI3d3jgLMUSQ83IBUL8t5Yiw4M7VE3BS
A6UzwYTJYTfe5UbGNynBNf6JBmu7efwW9tIsgSMrxIEpHs/g4C61Gdwb+B1xTAi3
ia3Y+Cue+hGD0uHRl/0qN8IXiMvSCX28xRtEZmUiPSOKbmY79zHLczqZvP+YmeS9
+eZ9yJl9lRyMnkdkM+13PRwFHOtafcXr0zxYbREuQA3kNi5DtGCK6iEl9PEvowyp
aBqk4rWj8NO7iPt6LEg5InHt2mEIya7fijfF4wpSq00zF0VC/Lxa2e2aN5DecZtD
GFEByqIpy7OIolbsTmjnWA6YlAzOIeOlqETURwwL2S6fFPB9buUu2sqR/pSw4ghO
M31o9WOdhWrQHY0Mx3eg/gZ9qK+lOUP7JHAIMxL17RLGPslwZlSQqjvC1cvGIlcO
O2OXLXHRNVLiJxwCCJo0Czwkmxj+b0urlJ2CMuLCX+q1mOErlyMDDwdiOUfID4GU
CpEWhMm9VuMolCN+EtSPZqZ960M/90H5OhddcPBRqpOaLG6mhCECvnbDrospJKuz
bBzGzqLvrGY6Ubq+UYfqigCTEs9nh1hCdH5wCN0feiD82th76lTqnhbYsffVGiwA
fPA82HxVAkovO+7t0o43pi88jU5Gt0HYHf/OyQNAPiRBy/6+4IGaq2pnXw+vA0me
RsMMXK3uqWGGcJaY4FrADhjZXWBSwO6ZuWdVJPHm0UHNA+KOv9a+DI5vuhW+bi+i
`protect END_PROTECTED
