`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S30QvY6uVem+2V3Fi+9204a0tdUiBoYqkpwD2B1xEsebsY8yf0LMZ0L9QDcd172A
xApTeP47PZ0NX+G30LV8szpK5c77fApvkX1ATnNQ4Y4oKfiFwTMKJwdhKim90OM9
be63kyvNLqY0artYOOLjxhg0KKmvmRS37nLqHntRAw9dzKXkHo3gwCs38+KkhR3A
bRasBqdLup/d6EREbltUj9sDVY7NWm6QH/OTK40oy6x3OdMmNFZ0SgKzj7B7FDmt
3vc+PfuZOulVEoYm3OZy7MWDBV5E5VFIgRdsx7mQcewxAeEmikUi6zRsCtX0YtuK
VdChep9CO3b8RRg7jnJp0+LHZ/+/d52ZUizcEc0a+LcQjVo/QAMQIytb3pcLOzg0
z7lNrkE+9K3EuGXkUd0ipdjMY1ZS7Jq87bJQW/2i2PeZXutsOO8W9KGr1I0RfO4h
5gyxBd4srUuSoT3RamoopJT2z5pg8Ezq3bFQMw5QewV/QHxZY6V3x4s9U6yXiXaF
tKxJ+cKYkpLcvPrnTQbx5u6cI/SwOs9rlDBnJXvnIURiBhRGVdiQTQXvbqusOuVV
xsXebC174g+JxX8hlVUplj/munDzwBUCJJd21WQ6vnGMFp8dKIscb6k7w7RuW60m
cLPatpgFDAjLPxOrwYWleQIQfAkA8r2aFGtPwmxgAk8+E7byJBWmCac6DXGi0Yzn
shTenbdeKcJ1kOfPkRLqm7rLbFqDuAIGGfp2jJ1B9BzFP9vHEU8gIQZJiT6v7QCJ
83ird3PVdQ0tXwhPCl4g/LG3sChDGV60ifTRVeH9DrRjtbbeQdUYlf2Iyp8tK7o/
KJz0MNgdV8HPCyYSrvtk9+d/1T514noLS0mHDGGGnaaWF17PvCh1MsVJ+3GmtjZq
V5wPM7aWBevSIh8r/+/0abkAFhWcAHs/nyccHig98/LXtKf0AKnGsrv+wzBOIDws
3QcpTdTkvoenm7uNRZ70S4w4nKym9b2VMw1iB3sCFQkla8YErX53HdrddWeBImBV
5B1sfj0FnoljgiYohkaos8CDVjOfDPxOlNJXY+Pcb3HwuLC4sXJFJ63e8xOqVOg/
4ZkPDjBYUCyeg5C1qgO54NUhZpMiPJJ3h2I0MFkLxqnhDdmLS5tM3lWWqXLogI3b
pxtZUhvhDWWljB5vs3ZDkc0+MI8azX/3oAjXtwu57UBj9XKSgQs8msaY517I8EfP
Z3/MvlXmF6W1Ae0X+KEoiHqLWsvrpRZoY2WSBmcGY2C1V3TIJZdsblsOK5SrQDCX
9zVGeD2EbWLw0J6yFB/ur4gNmsbV6kZrstO7x/G+FKVPdT4ThbiqPVLhfE30X8P2
Hpi4vVqu27rYoagraCTErLro0DgrtwJAyEHzsJ1NjasM199o9nRHhIQR9reORhL2
LmDsUz8gGLLSJS4jECTQvp4wv8ptp5KAc1obQ4ZIe8C45KrJJjp16S1JvJCcEFnP
7rKl3EpMDaB2FnvtW8demcQrNw+L+xRoGlTPA2I5+tZdE8/13EdONpJJOvC5tITy
gRrtzGksiuU0Qv+agRQJyNLvqHKPhCUFExxBxro5S20Ng2zg1lQzQu0t7jUFffnc
7+krfRi1nt4AAET+s1TCA8Sx7MMke4qk2Ow+pJIKB0ohpSJt6ofZP5vlJu8AggnD
/6Uwc4lFdo12qL2aX/sDdIDcD1fnnrajBd2mjvW5JQM/67A3xEYKevFaOpw1Inxd
uIVhghh2sHZKz0ezsLQNanSX88stAzQepck7Tg9NXN0UAOaRrA6TkIo/gbnVik31
ghh3bVLYi5sE9d9o9WUb8o+lWvWSwYGZbEAMGlUF2l0HDV5YD7OWzaK/tx6ylScL
6KazCuVPR31niJ3IzVGaQLjobQZscibQKYUGCFrksGGh305YMO0JyFkH60C8Wswi
f3H5Md0BKaxirwOhP7QmeC+Ek+An3OYT1iYDFQfFAsDAuWCoxuXDYtBZ8kYd80+S
DsmCuxibol7/F4ILAa9EVSuVYHbGPHcaLct18Sa32erFZd1IqK11ifmhG7a50OGP
B5eltOkNkwtmJ8nHVxysdbAgukQHZTeZKOKhVmNsgnXCbyFlPwS9mM+++IWFKyud
wUG+FnYEgUG7ADqKNF04/MjgSlD2RkU4ZICrwJr3clmwQBYR1n902HMktgeJ5mz3
J8q4TAyY872hbJkYQfnie/HhDQIfEcLIobeCoKw8wGKb8MjQhS6GRdNewiXPJNLR
ZCkGr/4gKAI/y4K1JyH2Fn9aSwm1253tGf1VYiYX/oSWKGlMYp5jdL6xbH7W/6Ve
ABr1LiR1VGfN4KK2QHEz/Pq32FfURI6+ZmQgUuop2XRpXZIyUfRSa//cN7YZ1uIE
A9ort3/sDlC3Ejs5CVxt4esuhnYsgEiTCD1F+ETADXbbp35gFbVac8MccAzlklGz
81k6YCNqYBUvBawNXRJm8bS8WMuWKBWVyRz7vROgD57ea1UrBtoMA2rlocQ6BOdO
gmJTAXEA1ETwQeBnZOcUNXTwxybVDoJx89+7sDAOkWlNUGVyf4ZJGFu4mVTCIIqF
7J2+Z1PbqNUTk1Tpdr3uPZmxPGDWimODg+6wWxG9nj+4gBT7zn1FRETAV2fX2bYW
ZLIxPmc4QHM/YyRyPn3wCk4A4EmgJc5/5dxKmziT/hEbYvve+29d0pc+yCAk839B
+JTxc20HC/GsglK4hIiNKHnfL4Mmu6Ri1dh1CosSVb7Lu9dgRKinBZSpgEWO5nDw
SsPWmDme4VE/1iHmCGfQZ2GkOHduxocrk3ddK5BtD+U3aVqumPJebDcG0OZomyR5
HmDDReR5c6PUxDpDHXyOuwUEJch+wLDm4Xo8cAd08Fbp+pV4lzBQp7mY2rE42wG9
6SPXZ+O9zc52sfcMuOrFjYPaXH0FZyoV3jGhAVct8iLXFeBTM0B5mazT/feI2Jnt
riuLeFx9x27HdR4TuhZ0Ug/VHEnFnf3YLIqIqb/5teuV6o2/HALypUxYO7GjqWC+
UvRmDn2MiMOk2Hos4gs+QLcN/qm4JHn3kdNiNHRCsCRkvwc6exf9NOrefLeWbqFY
zsydrtfyL0TgHI/Ur14m6iARglZh3V4VMnqPZEcQ6d0gKa8Nq3NR7NzIEqbcPFi2
enBamwSUxOoeyHArweZc6fCwa7CfGiKfPoD9jfkums9ej+CffWhWjdTUVdd3hgC6
F5qm9vPwGLfBQzw3IvkdDA/GqgtgyBfpC9hJPq8DkkAA6KU+5OrB9cWlLXGJdkuY
+o0w17nnN9Svib3L9Y2toc2LSGXn7sjNycYrrn3pTSVz6uPg4plxaXTX664RnBIU
Dor6JxwFz4H2Fox1jE+mnPNxNdmDSxNlDFWZs4rKWqKiZsRrs8aHV/oW6x2vEwZX
bRvJRKoFOJkoja4HnM8q8aABgHqjlgyJMGz9hhsN7BQ=
`protect END_PROTECTED
