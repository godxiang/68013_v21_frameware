`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOB/+iZ1nOa2OUXHc7DPRcc+hQljlDZay0MvIycnCeb2Vun/MVnyPjZm6TKFmE6c
22QrJZQ6JYn+dhbFrj3SoIqPmVrUsgMYKwu0LxGor6jC0D3GFZbAJg91wh2DnkqC
HtuOONd2RvMQkB9QHQCAyncGQ+S+vs+5x84ubpe8qeSC3u006JHUUG+hZfqr7MnV
/C16YURZL0i2xwKsZjRu9TAJv82MQ2z7U0ex1qLRb4uN0gN03wG7aP2pcxS553XE
eI3wJZ+i2rSAv6TpIYQXmwLCusdLHg/w6+TIHyZtnOTMJcQ1dYDD/Rw9RyFqJqfg
NGZ02zqwl2tlGWgNmZOdV7U4+I37WRJ8FZK/b8PJbPl++XRDTM0bDsEOCJDzUJbl
6t6sIvqBFR+6D1P2hgj7mFMJyk3Uby1gwF23WGo0w/Y68hucp/Ig8AW9q5vEONla
w6nSvCqw8JnE9a2Mb9088rWth4snzHTBYBfnhLH9I8uaWDykn3F12i7cTAcl+QQp
g82UCdeD2mGJ0UoA4ElsnJzvO41RQPyy+p9DWNE7q4G9OUFQeg05nAA2wYxm615B
4EA6to7EjuWGhOkY3FwK3cEAZpW/FWhGdJ5llivJ8f4Yy4jAZs6/te8LHSWQcFxZ
POKhJQRQBFa6lcjiCdwBzdvQPuifv0++Xsfg3MnuFd1YBYTs9e4bCmKHdG326eDH
1ngu4t3L9pT6mukSqR4i9iUu1uld3ZSACIxRpmmGTsYwUPfsDY02augC6z43rnF9
rZ1ebmzOks/ATVRj6qUtng3bydtIp3WjpFlgll6+DXDjkiJYAh2O1NY8W6s804p4
FwMpMzQX3pu0E50fxcv4iKu7yWEGrfCUlaKMhp4rX2yRFkZIdHO9fQBsChFakozj
/HJxoK/8e+y/MmtQy9/mydPaFdzBk35eAmMn8S3/8FsdJzj63JIhP+SmSut4Lqsr
9/SvDDfUGpsMz9MyPTqJV1EUM877gvCcDGalvBFEEgPjDMdFuyVBkIybBDxrNhx9
fK4vePfs1l07jSWmLhLmMLsgtLdf4khKExXmomtrgg/VJ6td9ZsSISlK2rwMwEuM
93SlD2n9futuFt2pAwz8dDcNLNRyQSFhZ9zXCaDM/3UaIpR4tGr0/bATqOcAepuV
HE2fQf2pTRcDYvAjah9VmObFiYyeSnedeXoT9CmZhjQcgCrxlJQbnWgqhMIdzfZp
0XHZ0bgsJPwoLwxkkPW/WMd6jKMTXWqMCNoZE1MiBqUF+ZmUj6xdt/zllCAI4fyF
I8xRDy88MQYKXrD18U8X1juuRQ7PpVvSA5WEocUYVu3sG1cofMMl/TuSzY/cJGa9
slZPisdwSoOiRgnTgdhFS2am0DiH+xmxjTXC8QZfGSAS5TWaa+qb/FERcrVwnRFV
qodRY/EDNaidTFZm3oNt2+rZyO7cnkbBZphy99LKkBKUNOVQMNqegDHlsLuL5z54
VTvluONc1GrObg4OP3YWFpO2TjHtn1vnWwdCJTdy19Hcgq7n8BHrD7FhWW9JafSr
5FmjahKBpgV0wAmzOytXYQ==
`protect END_PROTECTED
