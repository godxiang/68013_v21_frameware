`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYHFtqgWZy+o4StCajiX5FpN5YGnP1FZgR8ZhaQS3qRi3P/nvvaNaDNX1LLHRz8O
lBfhnSd3ivHK1OgF+YlEl1j20fjP+NDWVsa76ylVKlM8HiJNDuD9BurMDvM7ecqu
hpGnV1RAzElDG5CYr9zEZOqFSGYthm9ito8qRw0oILTol0WW2lOtJufoL6LRsIUR
spMsc9zzwlMDAZF3izOrX00T/odgB3RfVm3QabufMMUlmFaHeC83plVF6hR2EP8y
wzRb0J1Fgr5pqcQD3tC6dw73OjuhZ+xhmAd1LuPUalCnhvHvSNh8lyTkToLWyL8c
7IhZXwYpxMR9lsQG8MRsk4/l7mQ1BJ9yGf7454hQXQ2qzdPUiX2xhN8sMdPdlGV0
HYtUMxfWgdefQBtIc64ZUQUH9ANYApM5rexM5prCMI31a/8EBqCG5tXUZ+AbsE5h
ZlvuDKvTvnVgbw4/XWnR4izyY9QZjGuW6QDpKhZKkrGaRpIFVZpxxiOAUZJGNf1P
54Sll064MaDUL4hDjPNTtuwUPiRhwR9zaZRfXgqDjmCJ1d40KR2zTap6q++QVFJ8
R8x6mHLiGBMY799yrMyDli+GrWnPAsjteiDJae2yk7zTjJ/3Yqx31yWu2pn3erQR
qOwKv58CRjdNnFjw7Mp0CXbhsEQF/cx/OBLgC+2uGXraRhMHXy0bYZFp/dDhVBwJ
SCaUsHBk4OY/75FWO0qpIFatpFbKaqNTBGGVOLyNZ546wFLmNS1og27CTkEOOOrV
IClCRjYVPoo84mAQChxSITy8hssRAyHu049GpHanSnMXEkgk2nNEVH80lH/cwgkD
TDIUzqOpVBnN/6IiMB5kfa4d+miAiH5ISQ4JlXIg2Usr06b71266dnP+KbJMHfn/
tuuhIPaS4m9obar4fAK/6Wv1ixPVmrC9Jei6jFGwYlBAhOCbnN2fwjrJ3ZPdZxAt
Eto+GkMu8IuRwANWJE8HadM8ErfjtlvdQ9X1/ZQp71S0dHLFGF7q0tXjlQNe0F+J
izC2e9VeQcF0aFyU4OyBwlz0ehNjPS/6q9U3eDPz8qfKk5TAJMQoHtxltwabILn1
w4Y0hI0in9mjSaxI8juLpBalRW4yNWoNtKp+g5DI/6/bbHV5MCk7qHg9gNTl3G5i
BaLhy7OQO8C+kcuP/d1u+0eWBr+hmJ0MFRdzVUSmiDlWMKxxJaIrfioIMah6FK+L
DtbsoHJFvJspwoSrxbMV3iBsVIbjUjJkvf+5uHC2tNJX36l2v07pLZQLsnt5OYHQ
95VZrnoEddy9UdPKIdHg52j4+s5asM2KqAa+p4iqBWWwYX7cvmr6Hi5z5M2VlQlN
y+72sry3mf3UKH8NTxfVyVXp27BxNA/6VaS3SdgJTxnyv2ZrmBb48BR6oPN8BceJ
hkhvAoDDPqg7oYnJOSJJsf0nOnn2oluKYZW43agK1QcV+4aUtEcHhtFeEAX389f2
bqhMimxbgTj4/oxkYFOUTnfvepLENHnnXJzvtvJ+chyjEJHzTxr4LxdcfOE//COO
cVOPfHCDbCM+COSCUWKDip8Z7I2HHTo9v0ohzjljFiEId/wkVHAVcvzuCNUZWEg6
Bk9N/BOXfyBIhyelk1M0PHf764TACl5Tk+v0KJwzuvY2mrfVEZdag0jjIYsm35u1
uDlfKhdCDVZO516OWIO6y1yQs3uZpv9J/zziGqW4mkGb4V2Se+EpWtLO6blD7vmL
cxNjRsBKYY7Lc32+LxGYwEOAKzUj1cf/xKNhQ1SsRA4b6BMbhJJUdqz0Hti+LeIi
1PNYaQaXeNLOzATkSu10IU49x9AYTQfMTcK9CxLB2cCy38PBDNFSALpb50fgDwX/
0fl3uAMAJ+A42K7gSmacj2Q6V+fOHOQRugpmYO/1aXF2gxe5TVeuvY9vYsWsE4yk
2BWGVfQq2Ig+esjW7yP0AJB9YolLS/a40H+KyAsAL/UP2JQ7mVFNCKztdSBfo4l9
JRJ05qPdrlN1bWBHzqc3rrzkZzWOnH2LrWvWMGSpXmNNS8doa8vZlllJdkjuupmL
zsUsVMnLxMIEpauoV+8onJMCuUIQTYBIR6Vdagf40qrn0/GBruiTdF5DEr5lBvNd
N6PLleLJmUA3NVaqE1QyqqrmoV5H4iR0nACLdzu7/tufaOiXa3pgEQsFUhIYktey
MMHLzvnX7QxfKkwAEnk6z3TAQHjMxEQ0JzqDNDCbCBKKYdiwSghbCTxrmPIwiHP/
qEMrRXnsGfKyRmKTsBupW91bfwUPcbWZAhDyv6sTwqTLzbxquPY8PsOUZprAYlG4
h9UcxDTM5Bi7ENe+DNFO71rEYOtwXuS6iNXSxoZ/a7R+cX9HW5vNOrwlqRuYcq++
KAx0q98JE67KqpqxxWMrvq41ceXL89pbvQf5YzSOh9UkMhJymFihYYypRvK1MBFu
uk0MGBuNxGE+VJJqrV3wAhcgZ9z6WxRxSKAQYsWGk2tLzFQ9ioBg6r9sOsBv0tUK
hKzqc20z6ZdNfiLEaLP3IotPy/i9fHxu8D7UNiPMcktVof6NMEXJYyAGJQKaQ+If
oetkbB+LyVJOtK46sBlyDCAvB9KQHWdAH6ojpgz1MThXNT4zNQAvSfbd6pvKbs8+
sG4EILqTAx8kPjYoiZDBBdIJNJZG0sjXRuDjXnMACtyxbA8yw/pnpTvi3T3lhIGl
44sqFklSgNFxDJC4q+cC4mPT12Bw78c7de5mbakDc0mYVSO7NMcMgGouv62gzAcG
mkdNFWWtW4ELnI6Z6nR4eRDMo5wwQapSCSWGAk8KbKCfVTely1ryBe/yBBoBLPbe
9C/6YIc+NHyYO1HLTbRYWeDlcc0dJdnaqG5q2obC8fqjs8D006OhoAr98B9AYdg6
8pKU3jjDJwFE2RzI1X3dkiNOhXydtDsyJvUJg1Z8fJ7YD+A1NYF3kYBgdPkQOSTx
jHasTkK+xHToR9QLxpVfWBn65TFciJhZjx11v+uQTrlYNvJ8KWO/d76m4D+Fv/nq
VC7oFzwy18sR5TgtNkgWSNc9JM9iDn5k9bbfRG/ZWIjjdkyJeG3e1c3Vq/mp5q/k
IMHTmxqV73j9eQTUif7b9jdRblMYl5MI4rJqqJDd6PAqSsMT4hg160B6eEf8OH5P
uwbuS5FrEOqe6vuKtbVWpRNheg+pfue1CbT4lW1PXGnjGlJUvLkfxI5Qcy0BptFT
I8IHkNKBOWFQaySHj/c8C239tmX7Vsb6BT7me2aeh0nhJnsq3zm9sxUlIajkrLZy
4Qi0gHC2onwnK1QX1fSlqzlq9WGob+UlPcg8+iLhW31gSabte8D2M/9Tg/w4nwEQ
YL68qbiIvO9JFb4yeZ0TKANNvyIT+Iim75Iw7N+JJZiGXTJErVXmCT4yx9bIqdFA
7oW6kDNtnFp8TXija+V/CEvNr6dNGLIYKssggQ/XUR4qaaY712LWfFJaFiLoP4G/
inNLneBKj0/jV0iBIvxs6yObTBiAyHY1InXCNNoO1VOm5Kw7LpaAdajENOrX1qVr
D8pDouYZ9dnX3as25sjrWvQFR7+aPJUqQxCO9NxtYuZC7U6Wg0GDInGPgFnhuF1p
Hr2w5w8+nF4TJVRbrKLbBi92eOLVygnpDnFwGra5vQn1SCaQVDS4TxFXfuZUIGEi
TgnNFb2JdTLha3vkdlOH4EjO2iV/17L2/XYbKUA6cX1y/+uJMPt1rFqE79S3XI17
+QmXibIWNr5OjVkGbILBuWkPm/jL7un+YNHF+N8QQImC+0blqMhnKyfRB/fQuccZ
m27NpKP6/4ea1Wc0l0Hq9C84N2oYIdh/OUTXEpKRin3yRguxZj0jeWbo3A62Frs9
LM/eZyK2aRz75FYYtDsctoDoxiGGaA1HJQCn8YeWiEEDftdXNgQAUgvUQNSh4nqF
IStnmEvrM6ff+Rmr1ZRjfKJqDvRhrTq5raFb/IZin7JxqsbvUKz5dHw2wpoeGx07
PN0XpkfIjQ8wkXin9gI9bpNIOzWNMxXPghtfYX0/foHzx6DA4hjvD9k431V22hZh
6E1wY7qqyE6bM52Tr+FCzOk4L0LzSNh0+G3r4RnrTAQ23+Oc1HRtyLUIvnywqRPh
t6et8zCNR6A3npJtv5KOdduLe2yi+lML2ikYhgC0SfHKPs7XIHdcTmcgZ46WjEZq
PQuDQhHidT8pAmMZAlobNZ0pXzg6AZrMKare970/gchlu+tCgLwGIBCDw7wbBjmk
nYtPHs0aqP/JI/ty9v+7zlwzzO5GNbfPwUWx7I5cHMN764zgoePPUtAMpA9QyQ51
FAnhNf5I4Tr3wkPBFixWgPT7CNM51gHIinBWUUNBO3g7dHrJKVgYMFXRF3yNMgMr
RWz98vrDAiizF6/wU0ojqMw0vB07JM6fA3UcPbY2ZO4ctSyg/GNSwRKMRa405KMy
SvCjiFw6K8wcRlS3Cmmm8mJ5ZJ7CqXhvmjaaXVW9hUqMT2iDR6ufsHI4jdBA3R8o
i3IXKUfFcVKhA33TWNKWsr/GhQPzEiIjMd4V5p2w6cvEJmD2HjjcIK9rXTsclHVg
3z77f6Y9HMUg7MtJQKfDnxEzBe2nrNeRoYDS6N7xUld4TqWZV02mIS4S4Sn5mGDt
uDKwQckpjTD0zVVIkegGLDc9ILyxt8k4AZCKaCRbslrfrqmWDv8GxUHh3mLN7ujw
dq6Q4L512MW3D4VhEcM7/MM3zrZWmKQNtvvH5rgyI9AWZPWU76NxdtT5aIXc0GF1
hwmaZpn/rreEsZ+v8UQKd6fD1iebCVpt68zdVaiMDDn8kGfeA6dezchyd02aKnBU
kq6im/dXXhMLyMIOrsSnyYilnRvsMXKu7ox2L6t0w2zJJRdLCclns4mye1nAOI3s
9IwCRRlVMt2FJtER82PySkbC4XtnBm+xuQZ1Yg/WeZ1JoZH1DvWBvzuxqJcvoWy3
m7EoQ1la10x2fapMKTF1cA==
`protect END_PROTECTED
