`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3UH42By9i416PQU01HhjjHT2qnc7igW82pUiX6ScnVsQuqIj+947HOo2z1XUawm
hrRSdOxKmJnImf/fsjEldZv137+H9iVlBk5q/W8kkQXdxTXvLCt1FXvNswbnPN39
DrK3ZLtJNKBsJ2+otk9BltwT0c01Ycoby6Kkzj0/3sdWNQDyv3Rr/xf0EwtDqt9C
EYEPXlk5124DKrTs3zQazrIgwMiY+j55tPxlIy5YYgKdC3GZxCPI+43A3z+j+8cv
sPzBRINDnTHON4IuVFRETI2tfot8/v/jqFHI3A1/8Bj92EewMeuPsC9d+9YEPnxn
PKwa8F+Gx8iDkoA8dtywhfWkbl3CLXqV+T3tZBZnJr2QfF3/mEy+MQ4UmlUC1vsW
x10IEv9NE8Fp+fGOHgIZKaFQ0jxKXeMmxcMbCFPdhHzwxKspdkksue94/fR1KYxZ
I3Y9RHMJMuDJHcAR4fK0Rk4UpHMhlN6sIDXRag8e68nzHALbNSJJxIkbmJfEPAUH
IoD8SMVxLp4j/t40lMwW7XUAIPSPF9ymigRRi33AHC95o7ZSIzjJ3BBZvhiqiEUR
a7IsPtecqMVT7J2wzUvON9ZqL7m+/p3ljcF166NmArnjWO+VUZlt+h5lcaODEKH3
zny3dlWd7wjjlmLO5pI9rD4jwuPykg1TVM7uIl5xCfG117EO7dy+R0NThkNQ4jJa
bUx1gXh+ao4ZC0XXwIQa0jPa3TBAqZFwjTkhj3gIVsDfCwwcLiTRZXMCk9aF0YaB
/VG/OcHR+3CIqz7w/GzHt+N4RP81qkARJbfdxIN2nj2RUaDfdAvxOJF3tVdePfGb
yGJBe6CrnM4eoN+sKam4Mthsa0PFrtc08QxxUFBOIQ/ehl37dqf2PVFj1m8egnFV
J76Fy6e6DBZyFCnAdg+ga00SqNV4RdaI1l3jkeOP8MfGOafzANkhxmW3GHdjRi5a
pHLHIa9Ka++eymbmhrZgdaA0jSIDQIr7WDdfpdROMGX5reBRLmbmDYDReCYeuYMe
t5Pce1PMjGWhM331vIHrfxHBbEfQigNaqcP9raWYTsSogI72U1qGAjTvklqbnGo6
2Bu6m9mveOor6ji/zx8Cs4JnfURK4+e/5nZDCmgAyBlREahAWtN5zlSxHU/CFnhO
74KrmcJfG5jWrbshHPaIoFQ2+fXHwSwi4L991h8N/PWk/4EwvxQTULSmovtKNGxE
hoxyo0rI9e3E7HaHcGp1/L/g4OLMh9JOKGhnu0NHPCVghjPMNvwTCPia6h9iPCum
+SVBz/sVjLu6TurfoPzoP2RsI2dgtWQ1KCm98IX0uBTqD4dzQAn9Rdlh757uWrF1
zaxGEGuRaF/l8GNMOsJAn1EZYCbhSos6weU3ZGZ7kKwkATKcAhcsKMp8HQ/iZBJX
GxfUE5ZLdXSiNLEWpVD5zBeWIf2tZiAocRNf2Vsn/vyWLpgd4h7STFbn1OBbE+6d
KILsBTWKqNMlyQ3cHzwSu3iuWXhqSryLr/fNiPu92cFxxGEjR7O8yRx+CRMefIuA
WhyByukQZogmCnQof5tKtaDdbRzs6RIBsuhemRsBBpE=
`protect END_PROTECTED
