`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8GoNoWx+8JfqAZyeqwVAZidGW2W8LPdcqGPh0Vx1lqZsUPCH84ec9XmRetPVdC0
v1FchENoGEfJjg/1kmTfwS2NDkmgq5z3LbpJjfFfT2L+8zCfEZxCyK25loha/chQ
P7WDcKMwB0PqzDnqL13Kf/mTTqUFLaswzh7mtuWaDZQ7LKiYksIy40TNlwQ+v96F
dTnoMDtXPmfcqGXHmzOzYT8E+viHzTsg3UnsbpfINQYUF5xPW58mRnfqF1PW1NV8
Xs5MlD4nxQu8LWJ18bB37Yc5cdqXk/xF/2TKqtNhzsj2uLKuM5BAp6n9jNkNNQAu
PgJoNvtilpP0pd3aoCka/3o4Nu+DUHkcoXYdPJLnv7uRO1XQWoYWSxOl/7koefA7
CvEVXWs6ZI2z9os2Hd0MbvxHzV+p7oyvsROalCZbRZkfAOXwVinzyjHSn6K8tZBU
MeQ50akmvXzfVopNPlE2FLsmloC1+KFZw+fLPEjUA4/YC+OWrXoPxyZJYbxTyvrC
wymRGWti2TZ35tMcAuMiyspYjDpQKoGVY1HMrmU0in+wgMD83Lb1R2pU/pXLesZL
u26B1FbLeUs/nBCQg7GRb5Qn0fFiUqbhc2eoCkPObsxcvzgZY8u9V97F3xzQF8HT
eUvOLEXmmwio8nTy3iIB6YRM0vp9WCDwOqqV3lZgFz8/SNQ9ZwBr/Q304S6WJKMG
NEYi+wspevWwb4FqdJf2s2cAMB3Ss/IFXH4CYgneHnL7eG42HBU9/08gGJXSF87z
vUS6tk3q6fmtz5GPaK9cpzyvOtHCU2xKb8iz7IbZ+n4r2uICUeS4jxFBAJxzpEpI
fhROTcNDhNs/KjS3sSMlB9/s+m+eIj4g1+fEKbVK/9nr7sTxm2gmNXGVEe/8qr5i
iJc9LWgzFAmMqYqgDrH4QHVF+sOhcQF0yhPIS5uHGJO9sQmLCVQnDI+eQGAzgXmG
WEGLrONd7MWv3oOBPheebMT9cpI3CfvV7kYzPDoXpEjok/ra2mvqbO67wPlg34gU
VLPExASDAifh8IU7RvGf1BNGqLVFaIAhJ8Rh4dGP1eOna0kim7WQ/HKg3x7Euna7
pSlp800pxNVGvJIn596lfU5kc/HCeegdyd6WUtcZgrlDWNZRMbCcyt/1bCp3nkhH
FzKeDiRhANZukU7yCzLugUFw+I5kROUo27wQg4Ud8LtWI4VYEk4JsKxoMXJU1EiT
vCR9j9WKVgpOOyTU5HSvZpema3VkbUmhOHawJvhS6VmTiL81ruaAnlPhLfiPEvxZ
sFDN2wn1/aprFRongeMo7LF4+XeV36e4f+1X6BVHfEW11ZONrrr3e4C/BXeI10do
/WqLot+JqJtjMyQRVGPietYv3VqEZ56Fd7PGyUFp6Pmp2iqtjN+Goegtbg0D0f1N
NqyRzaBsWXsmRPcB/gxmfvK58e8ez3glIZ8ZruJRQrwFM2eqCZ2zu9SBA/K0y53t
3rfueo5rJXWl6f3+izDOMjfsDEuM95J/OelgwbFslph2aMOHbTf9WrI4hbtSN6Vm
+j8MGFCqOyXm1cTxi6MVH1hZP51tOuMNwXf9dSg3GkoIoeyYCQ5wVLcaSs1pvmlA
cDiZYpmnSekiIGIFu2eKSvdwNu+12z2b5wVd0unh9Xo8Z8EPCGle+1CWO2C6ueB4
ATVHc6t84DE75C3eBz5FTaqc53RBi5rWD9lKZejfUxs4vdL/2E/mQ70kaCcchaaG
xtinOc/08+7tqkhAW3HV3tCq8YgCsNDTdMCmY1h4GNLbRGv9erxvLL8cayEb8Amt
6VekUWM6e18Reqkl3cMTuPnCNxW05aVEhA8JnoAsYM7+7VH5TNmVPfwvemB7iSfo
ob/4hKqmn+sCcAM/JobkeDq2gvuuNvKhaVZ8kmQvlCIeU7BPdfy7Zmge5y8CNmU+
2eon/bHMElRNNTqpTJLhYTokqzxvVIMwRfDNCNaV2eGctPPMJo4mpv558t3zxqlp
I2iwSwn6RzPxr+lH4WYcCDFaRhQRwQ/jUemkB/VQGIOvyhg5HBNXlVv4jzch+tYd
d3EbOz3Pf5olWm3kGcCnfK54lmH4tHY6/qQQ+87l462KIAI9A5ai6xeF2+m4zWfB
Hn7kLz0vFk9NgvFJs3PicSZXrqeIOlZEeX30YO111JAEyo/7WPAfMRSbm23gMbbf
yd7eE00gbDCvNSuAfF3ABDiKruQ2RMiTdASpFIaGn9v+YYWmAmKM/keo63TYcHiH
Cef3wh20HRNirX1aw3bM1TLriyebbrBwC68QdkvW9WpeI3nZuJuoAkQrCGiB4gSp
0wmjHY8b61TFXUTK7KbSeJj+++MNOpI4rui1LQtJPYsnMHbK9FGikKzViHmEHLYO
tPsxpiaeKQR4JKwRjjGuZjjUDnRcO1TUnRKxcKUKMDZMkgU/AzhfJ4XEphbMZp6y
5J3o0XVfFARZAj3sWFFfWm/L1LDTyvhzJLnAE1j/BPojyQ2RxY7FdGjF2SylAqrL
WtfDDMPny/LzIlRKfegwgXqVwJyrl372SNPF6uJ6nFTpWEebqDQWocPEO8uDEVkZ
r393m7hG4MABnxIzgCmORyvUGb79DGBL0DepUPi54VhI1/OtP8xVJdxcoCAVGldn
UXWhaj0LlcPlwOD5WbvwBhkXOICIwICfFSfrF9fKOE9PmOmQeb75NqQMQckkQR8p
U7amo8cMO0fiCTDm8Gb5WBGUd3klHduFZcF1VsQtsEQbyVImowaAqVm798B63als
6ReKupT+k9dyzV8pHBsnP6CFEPc9I8NUXsVqSJgfG0p5XMtzrALug2rqpzUSaTKi
idTGSBmr+CxgbpZtgWD2Q7YUb3XygfALCt4oPsljX0NAy3EFiZ7xcadHZiBm/YKY
a7FlW69lalvgd2kSQBUPcLwyGKzMKYUU7R1WLbUrcka/BlWt4wyYiKP4hSNmaOol
zpV/StmAvHBV1VCvIPyT9b6AdsQ2P120GWNyP7UfO+YkTe9WpnccBroa5agj1RWH
flj5RwSVdmYJj4QYjqP1Z9cVLM0OwGBK7o5pfhatwYzI3K5v7qQyYoeP9KfXxblk
Rif5aIJ0n2CAh4S1ktBAEOMp+JOZ0Glz0w1KmDm5+OIB2lgbAHfS1eyU7dHziBpb
NG8VAdtKjw2vjb8PzVNScCpyRsc7skPZ8BcdZEMFzUkONhrNC4aoQ/k88GADPwSS
TC6icTehe0A0x4RLTfGfA9JCguU7hYP4JLN/yGWQmBu2n+B59vpN+HteFzCux1OE
msgTQWUTM++rgUjRSHRuB1FOQULAv/l0F5oMaCJeVvNArXkdT0Sz1xC+3idJ77Qt
7Kn6TJMRZKIUyJlz1EV//1eMwd9PUQ8ctzaznt2PDjtkDm7EJHhJ+sT3zesmbLgF
MpXSkv5Ex2AQ0hiVFdBRafibRhntoWQYZ3BZZiM+vZhLZghKV2IMVg44bZvPEMBE
JmjNeN+KkGou1EK2vGN49yUOqkf0TWjUHQGp6ra6lULQSJmAlDgHiu+12JC2Lo1k
TP+ImTFT3lAhpxhLhF2tHg20OfLhHwsDfJ/Mwk8qydOSBS+weEAO9IwVfcR/ziQK
YNONdgpjClLSbZhhEsWMd2YY1fjTT+b+8Ee4jHNrLYpD5n4WzDkhDEihCmLquhid
tz8aPi1XQXTfn59xAxyI6ZPnDBfl4mIWvV5zcQy4IPsuhN5J9bDZO/aiy07ErU58
fGFi/pY339ltmyG5Ej0FuR5xuxZbPzX83WrYssB4Gi8IpbN6GqWXjTLR1HXUzzrA
VzAwX6TL9twVDKc5aBCbD2v7Mzq/ScLsQHU+P7QHeP3lGAf6cNsut3jPz7lx2uD3
0dUtRennEZY0EcAHv1OFIyHnz1fxwXmxK3hUG+YwIbfFxKj62/M/Dzgqt+8CBiPU
ZCAW0nhJCdt/7pTi/N6SNYLwX1eidY4rg6NS4xxB2mxJjI6gNZXqEVvVf8GkDJ6o
OPvcH0msw8iE6fU8u35CtlvRZw3ZCYZo4DEKq0HzbtgcElTtMgWX1Wl7JbY1gD56
OVQy5ADDSM6wg0oqT7o9tibta6MvoS4yTNAy2N5QLlrL/qKwQSKZtW4PupaiBE3j
doZ03gEKjVHMOkEXv1oo2Bzbby7nd74G4F2vxLfo07Z7NtZ6KjBpgtozquSLuG4s
fHMxwuSe+qkK5TgvjsJgjKYA47VXrrE53eVP4HpQSAY9PTsKI2U++diF6y/FGW+6
2isC4WJ57AmmHqulMpMW9e+p45D0/i2Yf+LODEIgI5EtU6RqZuBOFZqVmhlXDgPY
AaxeuLn3M9Cf7AZXsXRlkwDoHOX3tiBUZk7n9aomUWwx9QBZDjkZvzoptTc/uAhv
RXNPQZO4G8j/glpoZfMngJUBHbDOitT4PiO2vKPks2y0wRsf50vQ6A6eze8gyDtY
ijLn8gtZTSWtHcthhrl/v1I8jMilx7C/nbNiprtQtyHzGdsNa+dkzyZKuv2cvLxI
Z2Ublbdn7RwHUmlNtqT1smofpj38UPGG9DK4a1OZ0ZLMWOxlFJAKPbdInYUGLyJV
dKcNmb83Vfj6vh8caJbb3UqLKpWca9d9dRRgxJJcbPNrSBKPWCGE134sSk3/W/rI
k0ZsFUNo20YvwpT66Ex2rBHrwuotMlThuNQfQqO1Yu5D2Wjm2AbyKtSeRpbofw0f
T/dKlvSwS0FxdfvHFoDQWIvvHXUQqWUI+opj5gzkOGZDMDJlLNfghwaog1d1Ahj1
639ggqUbBw+HnerImkDzg9wKqA/6DAmBselaf5/YzyZamZjk6YTTPMrHB2zHpKCm
U6cqylKbuQhrfCdvjERtexqByV7jLTy+IHudP/DDkP70NiprZ83k2s2zzoyxgd3p
SrUQaI1bdX7278+/BdPaN9goZ1FyfdECNkZiwMk3hotDycvnkKky/z1Wb9gtuO/M
wSMPzHJzTz+99SATqmIUh07z8Ksl7Hmzrx5ZNIqMYECXcmsfKO9KmY2hGtxvZqc6
+0cHEAu+2S7sLgumfVVjJYfHowRGxd0FY219ITrwJViFk/GKQ7Ey2r/gsvWD7mFf
PhykRkPrl/jF8WLVqSlEnpYwrTL8w4kP3a1Hi9wwJRbsJppgY1WNja9SvvUFSy+/
4IwrfmKWpFc+mDb72puwXRK6+D6HGuKTpF0haFEbRr9JMEJO4rDfUIapHHSmyeqo
2yvfgiHSCMAyXMFFY8VLuU5jqXUlF4EDAZtqPb6uHMIUffTn7t7huYN/olgq0p9S
JXNLcGeqYc39vTfaveflrdx369qff8cedhDv2bR4unTSZuj2MMBg8FpgNdp+2/ia
YvkCw7K1JYV5qETwLqMU81Nj1pDnfqspmXoHusrzD4QrLU6+g49xHgqFMwZ3z9UA
X8XZT5WygKA93iJ1W1DzAovhLK2AP/W7MZmcNFOccnQ+dc0URjmL50YRVeYmN+Hn
jbng6wI2XJZrAPrNvDNVtRD0ahQoFCkDmEqoY0+OMWgaeKm5wVaJCLQgPxhbxGl8
WZK/ixfhjywenfwGK8CcBI76KH9NbBVdA2iLCkeQNqNs54mleyGy2YExp6ViOov6
sotMEcIkx4Y9ykd158yvIUMefCb/BdRkkCmwZsDi4O2xAOF9zOdMj3yUHwx2uYLf
Pjy3lWvOHwOOSnGAWzyukiA77qFEqHkVZOcTlIwtmdPgg0oL6WqRdtdXgkHKO3Q7
fKXFlGScMtImDGXQpL9f6mbqp8Rt8VfLbfw4OdpSA6mv6fq+Lxpiszn1un0VF22S
YxVgqYCDQNhCbq4t0tI0IJWKPLfA4TCH4WCi0+aa+9wwa/4UvtemM+04abkHTq4Z
Qbs7pW1UIo+JtTvGQwaHAeH7SMKRfW04WZjBrcU2CBIdWPpwFdsF2s8EQW/HTXGH
Z6IVTDd1fFO/AbXPKUjUD58Cl7KAeDkje7Sx6nAFywgNtfwlDyFmcc1SuamKCrs5
kwo7RCugrBIXEiLkn+bzb3YeDgbFQ9yltKLpNaK1JkCn6E95dp3uqO/4QUyodX+4
5J+MzkyNc4SyWOlTGMgH9KUZhJtj2X8dNdih9nGqXFA1aTAW8YPrtOjoViESgal5
ID0OTU9cUnjzw1BpSX7Wwaok1XGm5EV3h34E5Jt9fnbdZHifIvFDqzwnfHoPtzB2
pchb8pCLkUGWIPSOQbV5706xChQLeFkYP64bIRn+MAp/40CLyaGAIPwGhGV7T7bz
N2sQzQAacSrsvWPMK6hKeBKZO1ERZoP9WU4a9ItpSAC0JQgD8OyuahAd3eyCMn8/
ijhZHbdAik8Xg/sFZ0oftPh1ePifwG7NbY7igBqa4xCMZ/lMyCcZ3aBOGWw7uEvK
KgJbe38B9KSQOWxob7ccAR45ua17hz65wiQHTKMqC0Lqq0r9glFlNnBfkRDYqZrw
YjWv13ITBVM3fNYqFx4FMe6isBk7s+25aLtvXxN0F63KvHh9P6RCyRAwUioVchU5
YkCBmVv6NeryMs4Ub3zUGmJnMUTilFZ3XaYxX4JvXiS5qg5ToBMW9hqK3nsqYuog
YvN5ORuPzqu1v4ZwwIjM6PeYq9osXQ8L1OknWTV6pWhg+bbIkO4+HPx7gYhNOUAz
p1JS1daIi8TW9g2A5nq7SQ3rkzeRrxPeoCaQ/7xW+xe9muo4+iRW0VBG+z0IRWos
tkGc1pNY5Zv+23ifQIxQdUThIwVnLqwGGJ1bvPZ6MEbPLSLw1c5iXZx4RvQzTLH/
d9J14LUuyMRpRK+wsX5Yj6IV6OQEVjcPKP2QOR1X2WPcjag3BYVRPY6NHCjBMnOo
mC+MqCHHCTDBsElsUAZw/ML4y6qw8zvjpoI/22xSGXvGPDENLp/QD/ZrXDH2szMk
MFLgy/XByhmxS4l54cG76NWhVqJH+1mizLBvAzD4fXeUHoxv/4NQRX0+KT/pJmGn
5ItF/Rvi7M9cdAHRlR1ZTC1n07OSsv/sD7q4YR2vVRnVYhVRXR/PIdYVBXB36LrL
sbbfUALUXwgW5Yh890fCRFy/BE6kywjxXn25euTLVHFJpJFgzI3CN9Cn2G/cvyJs
981TU+MOk5CZfOYffSv7MFw1KkJBSBCxgOqa2QkIegrRIo/7PMlanuGUYoAPKMpG
xivR5sCh+XilZXs01JSJMdwH3jzsZ5lsPlbu19l0PU1a7MmLNJcIpER8X/dU1xlP
G1Pr/w7vJxMHEilKkSpl+9MIFb5mwK8AoysrWOVWktjPwtaDqZU+8OQNGlRgEhjT
lfQ3KTgsWaEAi0o2LmsKR7Hmnbp2x0D1KoPaJCpL6aFZ0AP69XoqxcyEQLetHVOg
v6THAVbi7C5TmJl0m+Ti3JQKSaZM18TeEN4Qt5uQiw3vENBzjHqq2Nc+9m2E5JVy
5LWwuBXLKz2GurZ+CnRkolMTMAjHKvezcVWqWzbQZklFMZXsrgSKkD2vZnyXdCfP
Bag2Za3AZs69BMhMi45NV8sHjJc4ICkSRRd9+9dWiAAm/mwNdo+KY+PtDhmCKSD8
zd9JP8y/J6k/2ZH5KTTz1p0OLqvR0Jo21V7OAn9AZriFeva8Scdt5mPVZQlFHRiT
eLai7bhpD8Guk4zt++nqJts+9dBQy9cKXMXlh+SdmOFiSbssQKeaRJInZ0VFkuWV
LNZP3zOCpWaR3HnjQNk/xIpceoisSLJ7FxD2ircwRirovEmXQigxubqJjPm3qn9R
fw5NwG0WpRnvzV5+ZN5yIqlQFqOhdSWVdDFSnLkarPGML7RQrn8DBwfLGGcWDwRc
l1GxFClTDXx45Qa7rCib/uW6jDmtaVHbF0tFLy3jYI7IWO7Nn2w2vk7oiYnHpkeP
0nxqfqtUYmOlvQldF9+UqU8wnYM2lb3tPCkHVIQfJF2tzcGFzRkN/1EkXBxykrWm
KJcDGkzDm5iYkPgPyUZeTnm1QmLoo4DFaetngF8ERgsw4lNmejXHhm0tGJdOifdR
nKnxuBxYo99r3DoAeG/Y9yemmj6zfuF26xXwhBH97wk7KBrf1ul92FxWeC0SW5aZ
AvDu7S7vfF1WBS5YTCldncikyeBVJ/SnSCGMc/YKci/ehppJhEz15UwCv0B1yWID
pMjO6bZ07sp916fiiI2GIbX8A1WSGXg5Wl5t9DW6oIXosZ6mzyeV+DnZhTy9imu2
5kes1mNUfbzaihQgIQ+CrAX6S8Exd2vXPnZz3IAQU8fVo/L78ffS0JUi92R+6Jg8
dZRioTAmPzyoYXdgsz66CZd40Tg6XC+3ud5kisXvlY9eKtWQaA1FEPL/M+/Ue2BU
4uPZhwxyvLMtHqRXy8q0s37FCYGeRucG+qF83b5x8c/TOsf4HKywoqe5+lVelQ6S
Y3v5LI6D8w03gCsgbRxgAGjgBofMo6FbGGrujhnuq+352c06TiioAAf51x2hZ6vJ
sQNCxC+mZ9X3EFppGzINbCU2G/1toxoHS70vuxA1AAOPhxislS6XI6aI/3gnubhH
LU6IgOMdrk4dEBq+MY8Qr8ptNQt+LZhqeReKTxDZR5vetq87lQobn5nvrYWTy09L
CYX3AywxUWn9yZ7tRYcBPH6nhCRWigu7XT3tQUERibY1vLv6eLSmaJ2O9Xxg/cXH
xF/ca41xcYt3FvErXjRtN5v5lWDJvz7XFs+nkTe8MUlb1NDBLtekxj1WbqdvcZjm
olWZDT/+q/+CVLxaJd3ULKW8RUpHq6NB/94GeODWrLAt8d1VmQS0ormX2kmu6mcI
aB5tbxWpdd87p4mtg86PPIr7WIBz//ytRpYWjvEKeQ/3LdDeL2iQvdbe6HbTvQOO
UEAraJyuxWD6D+jmpCVzctwVNGsvYcAnLvBm3rVrS/75zAKhAt7X5FQXBNoJDD8o
htjZU9luBrXhVymQQwQDNcyB2bA5Mk7+nRTbBRKxq1kBvrJh+ck2gJMYRq4mmLiJ
Ifc0sftNOkGI9IU3fxhuQQIOQEBy82mY4D+D+tijWJMm0bLl+1NvrxKlYnYxn3vc
wOBm9RnzvpFma/Dfji3OLBh9I3TNPXvJG8aqb1Z9LAvU6FEiFn9xq88FNgwhn/7V
5Su0Oww0LAUeyVjGm5QMAszSvawmQp8hC2GnOVgmywQsVLWol9YPnvuZDKDDBrI/
9/eqYHfb+HSk5cJzcHIKUd4p2ZSXRb7chvqrGHFghvK01CkToyeEmTbKHVtDrxO2
A19ijGOmT5+xIFc3v6LE61ELTP2GAn3BAB+kJUEcS2dROxZ4DBlUxY9jrw6yPrZn
mLEwFM6k6NtQHJHBUAOHkn6jGA7a/4XmEZRINBrcDwRVvlORd2ledN6Y3oY9TciD
rWeWkgdUvPBgZfVPgM4gOs+kpYF0eyGQ8KLgbkg1fW/fPQcPcGDUFeRvG7/BXC1Z
7sbeXJBcRJxFdntFR7H2Aal41cyNW0iuFSlH5NeISfG7harjXay59e4efDT1fAtS
hHZ5gHT+s3h6va7JZSxTPkl8mAb0e2jdPbMX/Ry0rObGKW5htRqKVhGfvdwskETg
pPmkh4XL9DhM9Ukl04VorlUFfm4kB6x5LAAWTbv0V559Lp2EmQuBprayxmuIXqtk
L4a+9dnjeleFXfm2oKUQwvKg5ai12xKDeQ+d7KvwHJlhKk+6c3Iypmbk24CBcuhb
QxAOpdoFXKV8cz1hVx0XlacZq6p4SRo9EY6g1i4mFCE9IbXTrKeg7OzPvD5thHYC
dj6BMzQYasZZk32HuaCq6IxbZF9Y/yUU9gsDpmr71WYdtUFE4qX6LrWEpT59Bk5Y
xqe/KazqSHCBFOWPLbWesqd1+f8dcJLf/TUrngVzzET5yA0PLDwO+SKy7uPMrBNj
z3essfdGc8hUm+mFEWttN5qus9h7qZFsvJ4oy7yhhAZ9nVlH3ftfP7DKBW2/Edua
n4f8wG9kYYrby23dSsc5HidhJhLHKBWQVsQhSsgKULVGdAgUq+Ra1OM9ypI2e9PM
48Zg+0VR8Y9m2aO8bZ4Nwry2JKD3JXVg6DPWNkIs2Wy0+VrwGsRDFXZexB/4kqlB
zz9QHHn2UzUhPYRNZGUx9rOtyF0e9KVKgk1lXxTBGOMLvKmCEkO7SRvZt7Gr6Agp
Wdu+73qxJpRmK25FuOIbrasa/3xdj097gspKogzmUNKgAetD2qb6Jfuxildr/FZp
Zu8ZcvhV8+SSGdk1N8I0kdjqEdQa8DHrvLeY+ov4U1nsSFQ2ZwUuwOEJfcx4TIS9
fS9oZVmbC0U2oN7sAJZGKItue8a00lY/n6JO4d0bme4pA0PFeR0Bd6OhkW60Z1wt
d5MTMZSiP+P24OMWPsm62oXtki8lp4/eObIWbr0+OGwJfZ9kMCvo8hljZxjiCTxm
WnkGdpJJZYKir/byLOAam4OfGuWQ0OZE0DHo8yN8r6cIM3gHvrOdXfJAFCDiW8AA
yiRimkmvZ2jGqAeELJ22aJSvuiuX7sCN4IfeYcVgjt9FFtTDLsG3xwTNln4J0I47
l4s930ikRFWK+7wOjsP6miODE30nbZ7Kf6OB0TIkwhB6O9rLg8Egbw8GDNv0a0uL
x+sJKP2b8Y1BL/D1DlzZvXZspfCFOWDict6lq6DN/GiZPi8OrMGxI2j0kJxaTBJT
yEWhvYzbqYqt7zPrzaVkzG+RNqFkyAX4I7bTarM4id5AEzBGXiTv3LRSEnhMLAMJ
3an7qV2GIcpRfY4Gg/RsertBGut8n5bYQk8K1b0VEzBIPlxgvAFn8WN9juGfy6NF
wWiMDTy6CkiVTDs0ZD+XWzU9mfg+gQHzGijK+IdyLbyZKaZ+M1HrRP8p/3bOZtZ5
JgLDOKVv8ocfL1bzPabXUBkqEBfrQxOb2zg0jRCYy81OUVTR6JDDW/e+ullPewwQ
ILE0Hl2r4jGzo2elT6LIq471diMbx/2nRAmoRJ3MMfRh/7Qx4duicYpWTyX3g8Zo
S9IT9+JnTSEhyDMx9NheajvrrHCIziABqEo5sVg/E29eK+C+QrnWAVVLQBAG7y15
KLkkTgQTxbRKxYHp9iCg3lex3dlZwmoywyIRQDMhNBKUtT6Rm/o1yS7iWXflis4b
h5Dc/0t2DVZMbN7DkL/z9JsuPQC5JHYtH6fsYqyKdwoUUUmMQxaRAhwMlQKWGD59
lVpJvkuycADW0K6HoFm6JiuFwMpLcqB2JR+R0j5YHCJ7AJOvd+0gt+VS9iB7hurI
k903iQZXBMLbJ0rxLoIhK/HbxVjn+QXXH1eh7FBgCA97R90MlGRk1QQp1wsAMmk4
go1F1hUJrKzQoeng1SsLXOR736pEQ13+kgrsPVRRz4NoKLHOaKz7ltX7QCsjdZmh
DIqU7suXpEWVwXDdM3c/U3qF+h41IN0tg/f9GkBKb8kfnbRfEYPj69XxQTANlIBV
HJcXt+Ad92T734eApb6D8KMjeSkzzUfwUAD6iV0HnuXop4k6ybTOLU/KKn0T0Sxz
cVvn8O18tfbP7fEn4YKqAZNX2hY/ygAU5VxDQg9XfqIZXeM6jdeD24NqLeBOT0p0
ySyLuJUmX6U2aQYJN+bOM9wfRVHnBzmKKZU5f+t4giNGDfDCsU7a5r97jLfZQbaO
9V6Rx8E2sxFs5V1zUKLHUm2UCBqDo0pBKmvC+l2haAOVJ1MN6KiMzDapTEw5867R
Zzta64NnuOBpB6E8+kNL4ovXnwh79Eb5rwUOKNV0tGEt/ba84+vN3kXwUskmK5wy
vX4oJrBbkc71oA1YqTdfjcWQ0PX26O7Zlq/PtN6TwbLZnDa1Re7NyB2BIqPE47qK
hPaA5C9Q/q7e3ftzTS9t+CPU7CPIk3XDiJgmBVX9j6mGqUTX6UyGlKn3KJ1xvm1Z
pcZ0AUimYGPRWGkmQcn561hNfkBKdH2voW9x/Myv1MkDRQiLwUqCm6vdnKmYvgHu
7v61yKs7kPO2L/Nr8N/eQMYSc2fL5k7v/B2znRgMOR1W6sfSEN9LYEFdQa3E3QcO
LYlzbFWltJ03Pbdqp+gqp1kI+g9cFAKqy/LiKV8wncb0GtlcZX2fuE3vGJhdkyre
hvYlbDTo1EdbD8bzzmlvOlG5xoaqyepQYX36YCNV1xMmQBVZoT0Lz7FdicaQQ9Yz
D21Z3VW8XunAEs449OWDPza9lJSablKI6PntH4zc0P5fG6OVV/MGQZakBIir7k/y
1CGmF6gv67hXZzg5462mmtiqj4b8nu/2V0VFTXl4ksx2GX0xh5LqWAkB8KvtsoEy
YMX/oHoFNvllxqWXMXpZWhFMn0KjovQsq1rqA3cc+cP/fnFpoz4dzvFAXx+wCvqk
MDrPEx2b2q9SXKIw47QkXeN+8Ih8i346nUlI6XMnLSmhuwesfh4bavzgD/vKRqtg
x6PsuCytT5/KZo7TSiilH3RrY57KxJxqxr6Lemlo8RSAsL/k/FJOloZfgx3DT6MG
nZ/lTAf0LDkh2CibBTApHkfB+gVxFqLmTQLePwx/gvCTH+5QzFOvoivqGRcinIzs
D31ZlavhVfwSOg1Bw4/bRwu5eo7/3JhfXJoVUwCXqeDhd4ntz6ezrJXX0s9QeeW9
7SSl5Ylfo403OYlZFOQ4B7w7mWrmsV4p7F9X+YznVzRioZ9IINNQhUaXxP31EqGA
HIPDZJPBwJrY3LuhPUAXnhZrZI9Fid7BOgg7xbd85Ut5mYCekSXeyFLRhjT9AF/U
67RZs7Fix6NhaONVtzjFTZmgG91gB7t6zteufgaKwDfqC8ybNMYsiP1DCZuNvpZp
x9Ec/ooeajkJezQrBlgNYBefp20StJNloR1UI38gh5Sc+3RHE+Od2eNtFcxWRt8i
TiXKXEoI0nABrskhlOpHVt0HLAcLtfEcOQLEq4nafmglY8bqIkZzPkDWs7HvfSyG
DvCpEijAlNPKRIUUbEZWHwKreWFshqrxTGymfY2lh8sDBy3XLLpqcWDReKJf8SCT
7sXdHGFdATxjKkBPPaqrNAOt4XhUJi3jDhM/lxybVpA/+RE+epuEEr4opq0t4rV1
iCWWgKsdjp/XJVnkfHC7BfS9eqc3JEAQY4UtfM6UMU134u216q+Sj856Nnebj1Fc
ZtvVuyQl3lDCoYS/fAg2F1Lm5h5cSmNRXz6nN4Fa3B8ESCCmrrRu8o1rkiikIZYj
MrZoFZMizgshIt88uyhkWsPZC3WmtlrS46WLi2fIGwYUzLGg6ARrjvhyeQxHmWR0
wTk+80MXocMRDmoxlYnUMd7+oOKWYJ6xcVILGoucjDh5lsJDEyHZs12OaaFdLb7L
nJEAx6+eFbQ1HX2pyUJUOGDzaV3eijIiet5lTMAuqua+xPiMoYFeuNSV+T1Fcdoi
`protect END_PROTECTED
