`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhQPy2Gma1sSCS5Gjn9bdVFM+6LqWahhjn+MNNWoYL2CcJ3lPVby9fnkPqbmr4Yo
qGFO5rkx/cCTHZH1c3wZybvQkrntiQ/2inE7T1sPQIgilO8/v1PrezKxARu8IGci
OJ0RTiBJA+6Jd3auLzIXwvgysn9FiUFzdImMIEvabj6oTZGhpf+AP3ITOkTUknSl
UtoDbS4aguQlpQJ14lZVwHbDjA5NAeb2T+EgeKuuri8H/gtE9tL6UKC3QFfPUDW7
WC195HhLVsQA2zyOFYvK2wWphNBG/tVces0yAFz+tUsj95x1VIRcYYnXMnew+ivJ
mfNcQcjVadywEH8yFPVH0gOIMM9nHIGYgvcx0936NWgUgFQBQA/E8wQ876VWaJmY
6XrcPRdQA3WB6oQ/pVf/THyBmuG7grJCIedrHoXr9dgdGFBuuVUkaqb+WmApZDVY
5R0zvo+ZonpIyR7UxshYWrnpRJWY92ZnYbkLtncW6zp44gJU8rebKQ6l3Cq7of1W
RCdt2cCplbgk6zmROaZw7pmYQADIWpb2m/G6Ia+12TUKnUUI6OJczOhJdiihFPHp
k8ncYoV13OrnqqOIh0B+DNEX7cqtmCGKfFFniVRijQGx3/8gH8potmyuq7PwzJPs
i8e2r4Q+MTpU0Vtm3DTFo3Kaqi39O3HwG+yJycMeZlMxAL+4XrJnk6KOgcxqXIpk
zt8EOwBcMX+BEXa02BjTBk7ocf0qfzCd9rJwS5sZxN5mr+NCKBwATNr20O5VpddR
id5xHJo9aku3jH6XrSfpPCHuv6bZWT7oW86W1BX4d6B1OwrqtvOww+fBN419urdi
0gLl5IkWj7C+cXD3w56O/9D24GiuZ1TQVqd8smpUvvW8bvQuglC4WHCcdT12DqkK
zDRch073YWiKOTzSFILkbGHvOJdYjvXny29vt/3ryRDwKaP7Ibwe0xOYxeXJ2Qa2
7mK3VnR+5K9bVWW/r64E+oT3JfkdwHAkJNBnt24kEvL1UQHPcNGWdEBdrap3qMwZ
M11i0jqNUXQO0pepIWUgQA9EHmlvtoz2U8K6M9b6AZhO+BtPfTszpqaoES9ntlXP
DSEs/lumA5mNCPKib+fZFl4qYEwZ1dS3aMXzaIIgEV47fLQlk1wv9hKbobZl5Ffi
gRCkc+NXXeUoGnAiWWrBH4zvPbFXzrZePQX2/oWtOTKJh4SDA56BkjZUP7OlKMVW
9JNKojJC41XuwmaMF7evPVKHqRbgTICcKysGhkugcXWUswdEnmTUFLolvaxGmzEq
PCW+H78kGMYwjHEO+10liOSSrerSoYhbo1puqdw+9MBs4DAyRelKsjkJBQ0C9q2t
H6We1PesV7IdTYeOEM2YLmhk8udWwcajaSPOpBXg+Y41M+L+X90jnQK4dQ++QWW/
ydFAX9LC2RP2c9M813lVrsERAiKgmkYgKT/Ktrw0Eyn9GfLg2c5IKT7lkjemXwxc
6/Im4uIevd3dnRz/OQjd6DZfTBgZJlaq52if0X8TzhsBhDzkYsSP9T4XxJAGuPBo
kb29h5y+LTFrTQdtlFkWw4w0BiVo98vi2magJaURobulEIuOMSN/4lENpw6kUpVw
6NU24uA+3OkZF3KbM1KGGzoQnx7SV1WUK5NU+m9530UPO6RQiB5G/lnvyBOcyLX7
l0Lo2o9TABoLmoDNgvCzxu4d1sSRRzQP7gCf+l2KcG+YcgJvvlp3I6PJJ4tSqeX+
QVwG1aTxfPOtPo8j+xaLiEbgHXG6n5+hR+mpK7VMQ04ZSBfGtff6x9Gl8UfbEeU1
odvKjQo0UsRWesLMVqpuGk2Zy1fVUjhZ+lOI1V/Csizqc0LzObiKRE5JE1U/vDwl
OFgE+RSg0iUxVwyK4+QA7MY4dI/tU/4uKmUgCgvjXRB/u4YQtUJtngoldiAzQOkg
6Do2Fnx+iVh2zhKDsbYCcJVc2QKa6i+IDQ9U5zSPKpIe5BpmqARCxuiKsHbkJrJP
Bcog45mraGY2ddOs8v4VifI7k1N6xamsTJVwv5o+0WPFQvFybtpd++3OV2x/z0Ge
TrJfMeOP2vQ7mWcuNHCSnOWdcvG4TDBaDXeZnN4RYUzoEA5FTYCK4fGIQcrc7CBD
zcrahZ7PuqPo291mPZHIDKsa0OczZVyJqDwKchLZvl4=
`protect END_PROTECTED
