`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyN55x0KVJf8G2dm6mA1AbITSpe1wIU15BAApnUmGdHhhJdHOL8m+82Xs21TFOep
Sup+IKP6/3O1NFc5YBei455DGu9r1WMStPIcHVPwXBOrxM3y1x7Pq7iCoNaKjzuK
vEVQJ2dFmRdkgTvQuAKPTrGW/lGDBgRFOtK6c86CIk+wyZusAeG8PPssmgl+XlH4
PdZGR+zUDWCglccRP3Vagev7GYjXcpg0uMgejbq290JtKr1U8p1QS1srh+diXEtD
xCyUD642JtIXrqiGPZrJVnR10S3ScwpMtDVOUnuMVkt4HGcCgtCGp65W3d5ikttz
cm5IDNi6PI4h4vnfwrrgV8RtHrIDqy8Hg3+WgI1ibNTL8noJjrUgL0ZVBxDQuW1G
xjIH2r4jk5jNtTUz2c11k4rHedwwx0pFwnpjTzv5PTEr/aQAQ1VQAhAqKUp6Cz5A
YlSoI/z3L1F06zQy26JXIXz9XEJ15UO/pQH+RXEp4A3/4xQ8TICtbcWSRmdfX14n
sJBoWRuf2gc6wT2N2RDDspySeLuwsNOg3z/yf/FKr1l4+PwHqB4CcxOpIjgb/kEd
DDkkVFaL++lQoTwaY5W+w78/5awbJ8gV0jJpQjHfq+WbITe09nGw230nwyQb3muY
d2wMR6buw93yVd+EwJRlEe97lFwXyreUT/x5QFrb9m0X5d1nJRlBfA/+vTJEX0Sn
6tePQt9Lo16zTkwSfRNPDOnqTUgJY5aWZH9dTcOClYKtKZCW1p3OMrBQQUVgw2tX
QIKoaXRG+ToSJn3f0PsQOstONyMVqIDHmG103lUK3iLEBP1s2yUXkDJTQOUl+GXI
pI8d11ggJf4uMhe44r6ateCAWz2Im6fqzAd8v0XcrG7LDvXUcBLf6PsjkXno/Xik
VQ70NarJScCwqFVYW+ipagmy+mJk0su/oix57AmKhMeP+J9wEHO+6161jZ/AL/Dw
g/KvfoWoKx1rnUWe52M3HBTv9brMxwaCwKSZ+2O1hmjBzPgML6dVb8b5PPPDFjl1
EPqqqo0NkxliZN6QeZPTkJexMZwmqgVu+UT3kxhundmRM3/DWB9uZAl5Wq74Y+cX
LFX6xKwpb6H7K8G2OApZFHMmtcLC4JTdfgs5D9TCEXwSIy0PD7t0/QNOoZdu4ghl
8jgQh/CYaGumbT62a1NfkGc+XIM9P3TaqD9w7SPhaHdPmpGF4FpcR/P9TE7z0n0R
scTg2z+eBWLp3Bu8mLXfe4oQxO+m2rc0vH8xL7XL8ua8w9Up5JnztglbVjbDb93C
yf+081mUKf85Opn2O2vu9ferYyWDhaGbZZfTLI6R1thu0fCt7/rnSV8FAD3zTBu5
EpnXLVYUk0quWhMAwNKHCY5fBmQDiLQ+iAch3CgPvGDyGe/gDPpyAd/OC8GpqUGd
FpefIdfAWq64LDQDPNUDAoJDM4Vy+Gs17+xgpFwGRjzzvpDZuh/OzqN5wJigG0Uo
j1IitYOVC+rfHZa8IW5wR/K0VDC+on6szVveCGWsF1p4ftAHCmC6CUoEhiSI6pLL
jeCD/Py7hUExRXm9UKbh/OmBf6T0NeM86GU23XEm4z1IBGv1hifTPkaLpjCHVBPZ
xUKAic0Cby5IrF4AfVT6H0XpCB5LhwwHo3ORyCVJ8b5nyE8MJ5hw3ygFKlaC7wlH
LR5DPhPQwckCPIIflPcUD9gHskhNrMCZpnWG5MB1F9QAGOmHK83XWqmGDIPzXSI0
rNZylOyerAATkIxH5ekmbQk62nidwdaOc3lzOoBaaPnEElEN5DUprzEYBDxFLZDI
KRUbLCYSKnrJLXFHfghHhtNZs1YPYxq2WswVVvyYG/haYA2HGwyfSKKTUPtuVjRW
w/4yixy8nK2yw0KSPuRUxjX104NLzrsiDoNeb1fAsn81KdZL4kv6ZoNjZ7MdxjYW
6lNANG1YBCZuNAzUtxMXliKOHnTNRqdmGX9YknxP5eFiEIZ4QyYXlf4ytYGu/qDv
Q2fYDiIBJ077BdVryUX8k8aMpyB55mhbOXw41Y/F11yc7FjplNZVnmGZfskChleB
crwGqKqmCs6bKOG6NUZFCJdU6TY3qIEiEWYnh9TAyy+ZnurtFMexGEDUeOpTsVrd
pL7KhejkzpzD3q1z8Lb0zyhvMohNnOBNV05sJCP/4M8GVKA4/aMdkFOyCL3Amksu
6bs3y6xqDbHBzNMYfGztiAWxrIslS6c1NMxJe6I0oCvOZ9QM6zxvGb0PRDWE+uLA
KH2eYo+8vTofRegOOSkT6qib8FSggNySCRiQ44aVol0=
`protect END_PROTECTED
