`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUKq+8v0qh1YHDaoyUW2Q/4Eq1tB7w0HYC8u0TNoDNgmHeNyzvrW9I+fPB04JCc9
Mut0r/vFGk1B48q4poRGpbloIf5etbhZkqP3RM3XDy3XBY3NLB3bN99r/BD53qil
axXcc5JMRro49citn3XxFZP7uVYqL7gwZBzw7yDdsFuH8V0C9xu98fR3zNEuRvcW
5yfGNdsgCpeQPEZAcXDkm5VENAnYjHvQt8JxI12eHoZRDqBnTcsDur4BBBzLv6vW
Y++HIa+KghES9NoMschea1utmWalpog2sx+7X7FbvRH2vZZtwiRJVQQebRRDoDIM
waNirCdwN183/h9JVWqNbVpSZ93Bv0QJCkhVV9lJmmegT/zosV7FR6yb34X9gsdi
w1DF17Fz5QMYULt7bivYOHFtb5DDKVV2NjLBx/KRBCSC4ELEJudjVuPKrpg4aIaX
wHPrvpFV+GodCzUan67b6DPsA4Y9JbUO52+Dpj0FOP3NAakomZSEJjGteC7J2MIA
CjskMs7Em3x+iE3PYhsZ6+gbsbZqQZzWPxXBiDQg1B6paIGBBBDq8qdi1oDqNR6p
BhlmHVawESMG6YKDl/syn4KlnIftNhj4k9lSn+fvhYovBwgIVzVK8LagUCkfOpyy
5RpZQuumvz/9Ks0uKUFlf/fRUnHRQJDxsuAPzrDZeBxzQAm7cQQRFp2+x+Hkjq4W
utk34BqOAneSH4tTwfUTkgk41Lc/G0/CzMa4OcAFK7lPbA7pfpG4X+tSkAg2ot70
9gkYUWjvJu6mUtaK6l4RPedcf0bsD3dlPNluT73YWJST+/v3DnyG8awE/J+nIfMs
jtVMErriCxLnLiMXgsNDayIDmiDHs8ZRqj3ybTO86Asr6Ws5mj+KkQp3/wOKxBDm
bWdMA2Nuru0tMxUAyMVPpu7cASQwuXuDbpKofKpKfIXLMMNcQn3L4Vc/X1yAU+G+
nz6Bs3w1qaCS9+iDdeOlsEwdRLBXQ0UFtPSegCWSzHEgBgs5+uFIXC9LCvTea3js
7jnlRXF47RWNINpK3+8urFTDMM7H2x0ge7F9XGGiYR4BMT22P2f/YQ9W7AoEvnBx
LLJFumNssLHr5jPaqDC0p0LEaDkDAjmVOfcG+WDHljC+eFo7gGEEvnyet/fq03R2
X8L5zDP9iwpz8hQvuYkPvVurzGVMf12Sxc5A1dLW1v088LAwbZNYkGkvh8vVilfM
YYHKTTRbh51RzKsO7by10+SFwuLeq9QMO2jkSXfoJtrvv8G9xtNV+/X5IDauXnsV
puNaUIEdc0vUtFmOVaoRy4kL2EqGJZ3/3KaBNIWUZ8oIxKUHueAS3+zmSnR/eh97
dhA6QPYXsIIEQZ2R32xHUpwrSfQxjwsjA3GTrXS1YHN3DfPhoYAIVjkG/jgR57Y2
szMXzCT5SwYD/wMfJyyifisxy7sHkj00vunr+fMVgJqQbGmwH+I1ggTOhI8IAdv3
6grUw61YGjE3Ag9Vkp0xTZGLDWOeryURYGaeFPccFZiV52e2a9TR0tDs+icjeL/t
18cIBiSJkhX2sLHii7FOlvGtzMmKLPf7oIYi+WX8r3knmlgsr2eGlUBUhBuNGBa8
XbV65sDTHLwa9kKE9egWZQmVuuFGZNTOpszgwflL8eTIny3L1bR07TPY+ZDZkHKO
doueIGZP+8GHGz5e8k/WFSGNQjftk17GK6fd5dU9Y8MYgciBB/ODEro620iqEGPe
3Dd6sVZYepuX9SS7bQHtvdBK5sqmkVI4+7onlyWi/OvHRWC/L8fX5aLZaXtUlFrU
fMYzGbkgmAQW30P2aVBqmu/6CuZkvEXpRzC/GnH+JoG3x+ZdFys6Yo7xu0ihWO76
j7xtgR7qV9LncOPk2uOFv/i/MkFyEWaXOkpwjuxs63+Ua6MpLEkG2Y4ZVmwZorpf
vn1JNQ2SgUmWXVbr/1dMfBo20K3vhYjRMXl8GVzL7gCnPNGHgJXcndBz/QsTI9XN
A4ZSVYnpC9r1+yBfyB2Ls/k58qQqYspNCP43iST2S7tkNIskppPfG732AJTffUmX
XFW29A7Wotzypv8P4yIXDoa/ckRiOyi8haTSpx1g8D3eM3zyITUmWvMB96SG/kRI
fKoUdkaMqGr14ZJZ2+6PzwSixT1ayjpgk2E5kTy961F47yUIrTSNwwKG34mbzh44
s3550y94kgtSC2dh2yGusfp9Q1dUD7b97/UdtNn0KtsYRp1aa32DhFVrcppaiQ1i
dD/CvpD8Qj9dS33WQaYa7HCdD4IcDAFFWwA9fMR1hRhWpuS+eskbZ5F8r8gcLL4P
myoYc3q5lv5aR7fGXAC2sIX5nphrdmhxTXwTZuVBEbj+IIUfy4kEZiS9hydAnAPJ
f2Xyxho316j2pEkLhZhj83gIE4uEnNDh0x5iYIZ+ETMIC/DbABH89hs0ZdLIkjFY
OFGVih9kfO1WFCOGi50ljQFjrSpImn+czs1YLfzunQXvkhfqrdJ7BDlBW4cP489t
ZuwZSe1SugSpK9RDboGMsTRuM+1Hrj+TEKB0Y50jC8MsnHz0AyY5mMDfSG6OZqUz
wETvpzqV8VMQKXNv2tzaoo6jmbfPUq1EK09snJqOwd3jiE11km2XrrqeXSXGbolf
D5u27k+ArasghtX1tTwPAraGmsaicxE7s7SCq/QSCRJRwuBmoMHwIsY6JIUJiOf7
8g8p5EMHwE0nmbh0ITrZyKC+2NDS2eWI+y9/IvQcjRJLFE+XUrhU5QOCsfzgWYI0
EdYG2vfS+yW+MowOF8y2EmVqIhvgdgxxszmzkKfGzkuKg6h97aPHbNYiZ/NqCdfQ
2PCC2Ic5NdIQ2UIPuJwyJkskAo5sgebk+OMMtkY0FUd/UvMmFhi22OrSYs07Th2G
6UGUgXtlL73CrICDD7f4/wJnaNcaGu9kFPPjRwT+qlnAmpDy0Sujqpi9UxyUOhBH
Paw5/0L3V3Rq2m8esz03lOthITPnITVDePJTN8d6iUpH3WX1hPzmvJr/Ih0nD0F+
QYfHOqrc6f3/BzNq8Yzl9PRbI+2TYw6ea+8UUCImg0LCvHMuR+ZR42AaLb5mNDAv
ysfVk5Q3f9CfsWSJB4gEbdZ62+E+HuMuxa256+yhswmmC/uK1O1W/+RTvEpbebYK
3Tf2lAiue8QDiFWajndsCYYcu0wlF9OZrikYYvk/IWjPIHCAVdn5fogNhY1TI2J/
QHgE3HbSd1P5hlJwHMZSJm0615kOGI6/OfnN1JgYBgrAg4u0aBDJM9BM38CQSdf8
Q49BCNxWgTIwzYQjpck64c8sFscPGEOanLjv3z7cyMBE99ap0N0Zc1YuugPfM/of
La02vjucDBJB9VtUbkoBkRHtWesLlBWHrIIpPvdHqkJRlq0RGAIcH5eOKA8wcBB4
aEerlp9D94OmFRKTAmvXU9zn0ZLBDxEIJLOqEp/ORZU7a/BsAbj+cncSF3SbNVw2
7D4M3WfqcTWZWVsQz3P6cBinXnE7YXPvwsVMITlJET/kmPWl1mUTjSsleHrq8rnc
EqGRu8zeAAgnEdkwIGkA3R3JIbvwGcn6CMtpHgzEEncKCHTtVEV6oABaYevR0NK0
c1H9QU9awFMiDTt2R4ywN0khsKZsB0k73wmlOZRlPOWWL32XGy5eOQYpn0C/lmJ3
ByUGe08REazP2Xc7t1B3vY23abncB3EUKpk5iRrFxs8GI5xAv7MpWIOKuXwYukC1
0wMIpx6ONrCjKmyLVZNQdXprIzm69+Uh3qPRSjk8tfgx5Aac1ZcCUPsnNy3v5Mq/
D1Efye46aQY5AJYnw5xssv6Js4lJnvKBq7uZBqXV++1V69Y/OmHUM5oR4U86UDUT
xcvt8wf5TgVshdExF5gPnlrkDYAo+8OgtEM0C+VIDDPbHyzFlzJuyA0PhmpXcLyT
hCgR+11K5QM6VZTV1thLcvWkD/rNcbtvxEvNwjuEba8Uj4dBDal5eg6VD7VYPJE4
omtMy+WUNzsQ9QXeIrztI8fJQEb44bya56UOSFwQr8Pn76hl0xwhnTEd7CxDTMcl
AOwdq33Q+xMxesb+3dKvrS1TBN2qzlLPCGQAgHkbsc/X5LZw43eBxnl5aKdH807U
QbeSpggrvxkECAQ20fomKYMjtKvKFxrgzGaI7hpSNxj988N9o5+v4QePocha001r
XlIumnvwnv77AhJX7RHQ6ZRuS776tjO6MvHrNXWdWhN320ZBK1uh92UTINfq3YRA
oBUSp9JthzRLmMP0EzP9zUIS5DaxdN0U3eMlQFs/80KePy0zA53DDABeKdyTyRS5
wlBiOykQy9BiRvYWARTlskWRkEoTPRd2nIpTWrVjSOEGjAW4yn2pRfS/CVQxqd9n
tT6j+4D1feuBn7hkqWRg5lppZKBl0bixnToNsEw4X31gSYpryYD2NW3NXmRfwL29
+85LVwiK5IgXlqJn1P+21uJg4GRXDPQCqxIoV8+b4IxI8IydrQL1Y4xK/nx1m0YO
H1JMxv5X3WSxyxUVO2D0oIA/S/57uzpaGADEcRADydelX6HsontGkCa8jMcN1gua
d6MJcv2m3zpozLZI7P+VvNF1hdIgx0Ip4tv6gVYN4QY8VVxYam73yg8XyYY7otDG
RnTkvo9oQCYkTBlBnBRlhE3Bt0JZpLNgBGsZZpMEWpR6pOfwA0dURXrz9ooGzMfW
uh3fVBlzV6k+lC5wY6d7QTHrncQYSPlhjrRW7YNJ9RzgSgzmActebTtOcDck/S0K
Q33M/r/1h4ckMVbbt+mJ3DPtwH6s+K5ISCItI2aQ89+GyNLXrbzos6w20fthfWhL
zUJj0/bC681b7gmSM1zjktp1A8v1Ccp6Rk/ZWqiO2z/RNBS50yi0jp6kvCJKf2JY
3U92myIV3Eqkoese1pMMOmP23MlR+pQw6ZUfw40mBb7SUsJYGwjC5pDJd4zD4QQm
VJQ1jJDyuOOjg9VdvjjqGP6YlN90UdEznxQSKSYEAc+RnJCm2SJG54gt/XbX1sFg
vKjO0y4MVVZOaINoiRM0W7qD0Cbtf8Uh2kpxUvNY8ynLFlrbsg/trjjqbCBFK4FU
K8+KUY7satn7mw+IemeWUl5CY1YsYMmio/IqEGAViuyUhY84Kwf5mULmWrmBzsn/
FKKyJpZv+aM+WXj13DwnL46tn+L6fOH6YaXoCzrb9kPHlTeQUzmWol8o/169gQ7r
KFKJlaqFmA1JgakL66CVq9WtWE+UUYJ9tpsdTnJpnoHs29kWwAmiZt3ha41zYDrO
Nmf9Xv3dzXok3Sklic4z5ObvPSwjQJ9K3f1ebqtNbzUskukWu4zgJZcqu00Eh+Yz
/I+OiEbmM08aKuAlUhS0oF0xMkTA4f9rVO3nz0iYzwqPKILe/Lt+G+QKfaD+wjQc
AmbVT0GOIvMnpJk6nuCEUJIrFxxIePc2aqDOcn4D1nYgTFTSrArGNzz2xkFf6vIh
yAMBKrTYeFWdr0FQQMJ0FjCq0wtVINuDxL8h2nyXw7DGo07FT3L8uQ1nldNbqNOz
bEsQJLWA6qIPvW5590pwfXK/JfMZmlr7nCUibP8UYVF6i1n3PIhIwrnhlJKrt/7u
zgBwmyrnVxFSgswZFbIedZ/nfUSLMxZ0okGbRooW5/1sL7LW+tcekmt8p4lnAxOH
e++TPUY07g4GcvD6uCx7tnwHCC/yc9WSRzpBW4loDEedlqn8ij2Gy60boZoqOfBH
okYx9O1oy7HKV7fKlOs4upZcOSuCmUFxJ5nEPqaC46Zg+9Wqb2Ah2TcdSgWA1+rO
Lq1GaEZgve+C7ViPpwfBIVbZLeiWnIJQBzw5NM0mDQcZbhR1MULjW8vUsEy+Rz0w
YwzIJk1y6BGMCgYV6XQTz02KWAFyddqua/2MpsbA4n1BrRLskFJDWXKpjaJx/z96
tnxrF/bHWbJkFgKh1Jief45CH2rhlKCgQLcjWgSgMuwheBBHQb2hoSAnluEYyJcJ
7keuhphwkX2SMblV5Lzq4aWmqRcGI1WwovGby2BWXyJzkX5EW1JEa8ddF3/UQAF5
qf3x2elAjRSmfmB/EJecNRKDwrBSwZMN4hD7RBZS5yMrV057A3u8HWLhgSt3Q3L4
BQVzHwUbSib6T8K/ha/o3U7+ROx4HhglHJULTg+eybDqu1c3UFd3DmcoZtE3QUda
5XaWMevPnPxmf7MJwjbqhVs4GXlSAmEWOxTku34G2lXLsBKtZvzq2exUlXDRxxLe
dTm4Rj/XYKic0TXbdiUg9pQMHrw8IvsYRP9MV2RwxqPNhLVIb7Zwsgr04SjdwHEH
G+3zQ3sB1SaATGrPJ3GyfDE2MENVBp+KUPxvw2nMi/8OT4kDxqEgFOx2rCeUZ5Bv
7siJBAaAB6mup8fGDYcwTehXc5Uyopvon6fqUs+MR7AIOfVOyLMN1nENzpXI7ZEu
vuQbNPFJrhT4xmb4vpsFnXO97ZeK96JOOSx8dMPrbJ27XsHWIv8b+G9dEqBJfaEP
JmxlwtN1OOZ6XVvHAAjT09S3/a1tohgZe17CCjKcbJ8Cy1n36jHx8CKAXjmvdsyM
Z8tUUy/Nqkr5Y6C5z+Pl3OapzonJ9rrT/SJ97cDtcdAoMS9Xw9qMS6SELG/i2/3y
u9gUiQtveasHecAArvSY5cVsNPHqUaHnbBND2WoeeCxh0qFXv4qoA9W48eFPBOO0
R513OdYjYxSpLiK74R+XX5BnJU6JDANwP5fGZFt8eVL8DRbjHIcLIJ0KzQM6I/qc
3IDLxwOtBJMta+ty+Lh7m4wEJ98Vi10x3NROv7IddtutGr8a/vuzKfQ8oQjMzmib
VpW89W3peQ20KiPsZfvTpShdbeuk74kfPppjY0GDHkSaFexP+2+LFVtXnhhdewzx
F8JdplF8mykecW2/UvC3F9TBQnZy1lTb/G1eyOENPRM9z4ScrratYUrwVXycmnPp
vuYqEN0BWhDaLqOWEVAE2soB1jrj4BTMH1NFKsz5zxi1RLXHOtfvzXV9UbvkTEU3
+BilcnMAoKAQwx3k5UJ143zo6gV2dw8+IKgiO4PdGuqTH7kgcnRGjyQSr0qFbnlW
zPXgtdjXOQCetWxxFMHFS/0AyrFTqvudORKSxYl9+UCszLvxiElTYrEV7vTM4GHh
uco/GU7EJT/TBwKDYLNVVqZAiwL03ELJEuSeuu9aMfm45a/9wO23L40Nx256kZn5
cD6F1BZvCBGq9RmbmVr0x/pWjg8uuNmOqzUZSiM2ZZYg+GtNEv1U0vAAkp4HRKye
XJ2I3p2K85IYA0Myz5oIk8xy3uLT9DppiLSIXghbLTH2AgIcdYCsFHvyo3us2FX9
0P5Fo7YjL76U9LkSIX+LysS8LEdzMcGtjcVlxP0nAr6W/wqW9DjVALpVoQ2YYBSb
Gqd6ZVn1m2aqT2ba7CCBo2xorOqeWxbisHdqqI3m/Fni/7u0MNtptnLVJl1s0WbY
n+1wcI8L2QYqDUNN8QVEYVavQxovlwOX/OA5VUulAg6zh7YX883iB3DRJwwcoG8T
qCh2H/QUFY+wbG8Y94BGRP4gQ+7MoHPOBkVU1hHjeTM9uAWJePWluCYPa3zH75Pj
1nAFxoKS4+wgGnuIXIaZg9+FOxqwHXkhw5aIsr35fenPzmp3kqoARcNq3xmm+em6
BetCg/NLs6Yk4f6jLbV6v7aBmQCoB5s5/Qq0ZX6Beq8OzBVpcol2q9lPTegrS4eE
zVoccKjrzp3/KLE4E+rbbFsaOWgdmJ1mKk/eFYS2EYYPHy6XzH2xOAirhmLFxGiV
okLQPtrZUWtUODe8DS0hlvnCUpXFZqTLSgzxXxuVhSA+DDdzA8rFVldY7CgAP9/z
IL1pZcciayhOlw1svFUgs9hyMbM7Q2RpA02aGneWXnadWCAyJQTFml6WsDPQP7nn
dAVEZs0fK6a7QsJvzjkUpPAZ4+/lVpHt+5QBeOTqt+jVm2ulYlRzmkOfTY4iVf5b
OO5GV4P/Nx5yjf8ErpfD8AWlme9ddKVkT86xn/gTjDG//gmNLPScpmIppemxIy4N
N3PI58q3OINih+ar8G2N4BMT9IlZu901gosBv/4aeFhg73qa0SFDX+eyMdPm1mv2
MYSpIQzTbLTV0fEYcJME1E8eRmg2DvdoNskcFOwFn6qcD+wYC2Udyilky7uXQHLE
zwawiWqVmcbZKXueaIOP0+OE+JgrtHijWsxhhUmCCoLEshXkGQAss7KDUSyZCL0t
H5cD/EPRhX1xyyxkbZQmx2V2OXjNLUiUfgot8egtz66pvGopnQxGVqZ3FCK9L93R
01bxlHmJXBemlYK2bqkh8NYFodqtJeRpgGpnytudsSvo4IhTlW40HDdoh/+Yt268
ExhmZEnFzzE6fvqmTWy1R1TRJjT8+h05TRorGKqPiiWVebmoZdFNF0ThjcpYrG6e
c3VMbGoK4drqgYFgUkHDk6q/njM+WBgqZZ1L6/NpRsnLkZVROWf6ST/MFYiBkwwo
rJAlfmINYnLCBvdK13ZxFmkasDddRzGRssKAkxOHU2zZF6ruKDH+5qOP1WGCaR3z
RjS6E8RG1GrTuX5fOctcVpn9RzX5eikzkwSkRdmWXrDLvYgaXfJCIez5G8yVJPCN
L3+mdjlK9cUnnEm6M446sdS4lEJSTqFx0c2sZBNXY7Y8jyfutr89aXUT14mLYy67
h9XpDGI9uHFvrT0ea8j/Syj3Ic50V82KZ9aomFB1T/f/tIqrkln6n0y72oeDZifE
BFwCbNWjIG8/anIg2HLoJM6Y0SoKs97RYMp7mDS7M/w7ebYFUEfwyCUpcLgjwAo8
/TUWrx2ZDratUakcJHgaOprEMbRhQ5a5h4eCt1KVkxQeJXUAKMSGp356DFCf9l10
QGyKZZ7g4h8mZmmdmoamhlj5ED4060E/BLZ/EojsfDOQniPn3DtFwRHJRNagn6wy
UO0ZfhHWq9gnOEKfw/W7r58bSVGGZ43qdppYtI9d8JE8Hr9Kr9KngotNjVWAUtVm
A7W0pRQtEx/wencoHPcoEzttSBMV1vgvc0odynghboMEICr2gnyhPH6WymMQRNRj
If34TkFTYG71mscUrjNLsAE4lqt/pYMuzF2+BRRNOBLS7RgZy1UZqJ5uMPKA9SG/
jpBpf5M/pNU3b+WMCefrStwA7ryBHS9Dz55FJDHPt2I36Si55yCQw58wAQsnY9B7
CREdxjBVFGE2CiLcxRD/GDtLK1XGPubutnW57/vVXKa/DKIJ1E3r9uM8T0OSnhfh
LvPmXKK6xRvRAZ9W4l3LnBlA/3cpORDsLsUUBCl4XWIIHF02lQHRrmjDcMB36UcR
CJ+McAM2tikxvP0klAKCGvYWX+mgmzbPcNj9SCOFKmU4P8OET7WqKuat51mChJRF
Mlk3l4SyUpq5qz9d3900lhftY4Czc31dQFCdpqP7KOtnxc1uYBiH+Is2mofABoGd
Ji7RVBTKjhQ26QVJGNzGqmihDVEfimhm1t89K75vWmmcHeT6i04ehqOPoJia4zVf
FIiHc5D3zWdv+h9f2Rxs/YnoOvChjCK8orCukfCqOrfUFjXgIuqGinKSXBWS4ztv
eL6HByduNkXUuyRiVUqyyqUxeIItExfNy+aw0awYxCYB5KQICcLQccRm/Pcbrmfj
OR9hvRgScmTm6yQRefrtRlnzywsq5szsBxxrcmqbbFb3VSNiQsVje2pUthwzgKzF
jbMadr7oH0hN7EnX23D/Xith34kHsVSv4UJfeXb57bheaYkrnch6PWUEb49uD54R
U/p3UTfLO2wYTmyda2Zx2K0t0wbQ1sEWO1Onn+QAd1aWBGXyJgWyvSgza+M9PLso
qgl8ILA7tDrDaek2ADe0VstogO/+1hBmbBs9Fo8i/dFZUQaVpPQnfySqcFWEf6qw
v2xTTj0ZZDUjyC4GOwey53SAFZscvWXDIoFQwtO3IxBAZnBk0OQIAfUB0HGT87IF
j01xsUVAb59qwudebOHtMb80nS/jgErKvYXeZ+jjoYAAdnYEjxHDqPDdSx3XOiYA
0y7Wa5Ms6ib2HB5y/Y5ik4+gH9wGFRBq42cmLylybJKKOCxUTrTk0OT96hXYcPes
FciD1hdqmHshIVy06UpfQ3aGWrhd2Wb8nuYEL5RL6CWWWn6ThTHJFuT2lwAQI3+r
OajWfKPOKb4pSn9nDDAfWdnaswZxwW519FfQ0gpDPq2XXf38R9KDtFTcpgJJBQhO
b1x6GUHUzGJlaRMe4gok3gEcnzGzjO7Qq5F1FsmLJAocHvB6y1t9koL2aHson72b
+PvSioxxc/xBibh8ValKvbj60phA164Q54fKM+N4owN2dgzyGEZoLbQFoNMa8xbM
Vf3BMWj1/p8a7VlhYp5WLFvnuTdWWFDH0KR3qCqLPAWpdR3xZqfdnAuB5cO0KP3J
fFzNBfhZnb5iGfkMFLLUod5/jeNp4mQuJy2BdQCZfhc/0k4oI7cj9Cz2xg6uoxlF
SLAd3bULXrZC2lqlQO8zr3M1yE+4zL0Pxi/TYsiJ2PWCl1kHfVIWrooSxzwplmOL
hz6nBsq6Yb2NemlwHTG6kKwfSZkAdCSeS7wytf22vkWgF61aPnauG4Aa4vgbyut9
tWcfQpxFb6mX6VZxLUwEEMyplCASGYNMWjB0d263UPzKoXEalWqX4/GTsB4rRUTE
RmFuRQcJWhGPjCb5Z0en24nghqprv1T1tqo+F/s+INnWzkbpKv2QnQHAKl9bMKGF
Zh7fhQmckFBNn/EYAeWkmGy22i+/pQXtck6giNRoHrw=
`protect END_PROTECTED
